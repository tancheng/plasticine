
module SNPS_CLOCK_GATE_HIGH_FF_1_4_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FF_1_4_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FF_1_4_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module Plasticine ( clk, reset, io_config_enable, io_command, io_status );
  input clk, reset, io_config_enable, io_command;
  output io_status;
  wire   controlBox_N6, controlBox_commandReg,
         cu1_counterChain_io_data_0_out_0_, cu1_counterChain_io_data_0_out_1_,
         cu1_counterChain_io_data_0_out_2_, cu1_counterChain_io_data_1_out_0_,
         cu1_counterChain_io_data_1_out_1_, cu1_counterChain_io_data_1_out_2_,
         cu0_counterChain_io_data_0_out_0_, cu0_counterChain_io_data_0_out_1_,
         cu0_counterChain_io_data_0_out_2_, cu0_counterChain_io_data_1_out_0_,
         cu0_counterChain_io_data_1_out_1_, cu0_counterChain_io_data_1_out_2_,
         cu0_T21_0_, cu1_mem1_N30, cu1_mem1_N29, cu1_mem1_N27, cu1_mem1_N25,
         cu1_mem1_N24, cu1_mem1_N23, cu1_mem1_N22, cu1_mem1_N21, cu1_mem1_N20,
         cu1_mem1_N19, cu1_mem1_N18, cu1_mem1_N17, cu1_mem1_N16, cu1_mem1_N15,
         cu1_RegisterBlock_1_FF_1_io_data_out_0_,
         cu1_RegisterBlock_1_FF_1_io_data_out_1_,
         cu1_RegisterBlock_1_FF_1_io_data_out_2_,
         cu1_RegisterBlock_1_FF_1_io_data_out_3_,
         cu1_RegisterBlock_1_FF_1_io_data_out_4_,
         cu1_RegisterBlock_1_FF_1_io_data_out_5_,
         cu1_RegisterBlock_1_FF_1_io_data_out_6_,
         cu1_RegisterBlock_1_FF_1_io_data_out_7_,
         cu1_RegisterBlock_1_FF_io_data_out_0_,
         cu1_RegisterBlock_1_FF_io_data_out_1_,
         cu1_RegisterBlock_1_FF_io_data_out_2_,
         cu1_RegisterBlock_1_FF_io_data_out_3_,
         cu1_RegisterBlock_1_FF_io_data_out_4_,
         cu1_RegisterBlock_1_FF_io_data_out_5_,
         cu1_RegisterBlock_1_FF_io_data_out_6_,
         cu1_RegisterBlock_FF_io_data_out_0_,
         cu1_RegisterBlock_FF_io_data_out_1_,
         cu1_RegisterBlock_FF_io_data_out_2_,
         cu1_RegisterBlock_FF_io_data_out_3_,
         cu1_RegisterBlock_FF_io_data_out_5_,
         cu1_RegisterBlock_FF_io_data_out_6_, cu0_mem0_N30, cu0_mem0_N29,
         cu0_mem0_N27, cu0_mem0_N25, cu0_mem0_N24, cu0_mem0_N23, cu0_mem0_N22,
         cu0_mem0_N21, cu0_mem0_N20, cu0_mem0_N19, cu0_mem0_N18, cu0_mem0_N17,
         cu0_mem0_N16, cu0_mem0_N15, cu0_mem1_net3732, cu0_mem1_net3727,
         cu0_mem1_net3722, cu0_mem1_net3717, cu0_mem1_net3712,
         cu0_mem1_net3707, cu0_mem1_net3702, cu0_mem1_net3697,
         cu0_mem1_net3692, cu0_mem1_net3687, cu0_mem1_net3682,
         cu0_mem1_net3672, cu0_mem1_net3662, cu0_mem1_net3656,
         cu0_RegisterBlock_FF_io_data_out_0_,
         cu0_RegisterBlock_FF_io_data_out_1_,
         cu0_RegisterBlock_FF_io_data_out_2_,
         cu0_RegisterBlock_FF_io_data_out_3_,
         cu0_RegisterBlock_FF_io_data_out_4_,
         cu0_RegisterBlock_FF_io_data_out_5_,
         cu0_RegisterBlock_FF_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_0_,
         cu0_RegisterBlock_1_FF_1_io_data_out_1_,
         cu0_RegisterBlock_1_FF_1_io_data_out_2_,
         cu0_RegisterBlock_1_FF_1_io_data_out_3_,
         cu0_RegisterBlock_1_FF_1_io_data_out_4_,
         cu0_RegisterBlock_1_FF_1_io_data_out_5_,
         cu0_RegisterBlock_1_FF_1_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_7_,
         cu0_RegisterBlock_1_FF_io_data_out_0_,
         cu0_RegisterBlock_1_FF_io_data_out_1_,
         cu0_RegisterBlock_1_FF_io_data_out_2_,
         cu0_RegisterBlock_1_FF_io_data_out_3_,
         cu0_RegisterBlock_1_FF_io_data_out_4_,
         cu0_RegisterBlock_1_FF_io_data_out_5_,
         cu0_RegisterBlock_1_FF_io_data_out_6_, cu1_mem0_net3732,
         cu1_mem0_net3727, cu1_mem0_net3722, cu1_mem0_net3717,
         cu1_mem0_net3712, cu1_mem0_net3707, cu1_mem0_net3702,
         cu1_mem0_net3697, cu1_mem0_net3692, cu1_mem0_net3687,
         cu1_mem0_net3682, cu1_mem0_net3672, cu1_mem0_net3662,
         cu1_mem0_net3656, cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_incXbar_net3602, cu0_controlBlock_incXbar_net3599,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu0_RegisterBlock_FF_1_net3515, cu0_RegisterBlock_FF_1_net3512,
         cu0_RegisterBlock_FF_1_net3509, cu0_RegisterBlock_FF_1_net3506,
         cu0_RegisterBlock_FF_1_net3503, cu0_RegisterBlock_FF_1_net3500,
         cu0_RegisterBlock_FF_1_net3497, cu0_RegisterBlock_FF_1_net3494,
         cu0_RegisterBlock_FF_3_net3515, cu0_RegisterBlock_FF_3_net3512,
         cu0_RegisterBlock_FF_3_net3509, cu0_RegisterBlock_FF_3_net3506,
         cu0_RegisterBlock_FF_3_net3503, cu0_RegisterBlock_FF_3_net3500,
         cu0_RegisterBlock_1_FF_1_net3518, cu0_RegisterBlock_1_FF_1_net3515,
         cu0_RegisterBlock_1_FF_1_net3512, cu0_RegisterBlock_1_FF_1_net3509,
         cu0_RegisterBlock_1_FF_1_net3506, cu0_RegisterBlock_1_FF_1_net3503,
         cu0_RegisterBlock_1_FF_1_net3500, cu0_RegisterBlock_1_FF_1_net3497,
         cu0_RegisterBlock_1_FF_1_net3494, cu0_RegisterBlock_1_FF_1_net3491,
         cu1_counterChain_CounterRC_config__stride_0_,
         cu1_RegisterBlock_FF_1_net3515, cu1_RegisterBlock_FF_1_net3512,
         cu1_RegisterBlock_FF_1_net3509, cu1_RegisterBlock_FF_1_net3506,
         cu1_RegisterBlock_FF_1_net3503, cu1_RegisterBlock_FF_1_net3500,
         cu1_RegisterBlock_FF_1_net3497, cu1_RegisterBlock_FF_3_net3515,
         cu1_RegisterBlock_FF_3_net3512, cu1_RegisterBlock_FF_3_net3509,
         cu1_RegisterBlock_FF_3_net3506, cu1_RegisterBlock_FF_3_net3503,
         cu1_RegisterBlock_FF_3_net3500, cu1_RegisterBlock_1_FF_1_net3518,
         cu1_RegisterBlock_1_FF_1_net3515, cu1_RegisterBlock_1_FF_1_net3512,
         cu1_RegisterBlock_1_FF_1_net3509, cu1_RegisterBlock_1_FF_1_net3506,
         cu1_RegisterBlock_1_FF_1_net3503, cu1_RegisterBlock_1_FF_1_net3500,
         cu1_RegisterBlock_1_FF_1_net3497, cu1_RegisterBlock_1_FF_1_net3494,
         cu1_RegisterBlock_1_FF_1_net3491,
         cu1_controlBlock_UpDownCtr_1_reg__net3581,
         cu1_controlBlock_UpDownCtr_1_reg__net3578,
         cu1_controlBlock_UpDownCtr_1_reg__net3575,
         cu1_controlBlock_UpDownCtr_1_reg__net3572,
         cu0_controlBlock_UpDownCtr_reg__net3581,
         cu0_controlBlock_UpDownCtr_reg__net3578,
         cu0_controlBlock_UpDownCtr_reg__net3575,
         cu0_controlBlock_UpDownCtr_reg__net3572,
         cu0_controlBlock_UpDownCtr_1_reg__net3581,
         cu0_controlBlock_UpDownCtr_1_reg__net3578,
         cu0_controlBlock_UpDownCtr_1_reg__net3575,
         cu0_controlBlock_UpDownCtr_1_reg__net3572,
         cu1_controlBlock_UpDownCtr_reg__net3581,
         cu1_controlBlock_UpDownCtr_reg__net3578,
         cu1_controlBlock_UpDownCtr_reg__net3575,
         cu1_controlBlock_UpDownCtr_reg__net3572,
         cu0_counterChain_CounterRC_counter_reg__net3515,
         cu0_counterChain_CounterRC_counter_reg__net3512,
         cu0_counterChain_CounterRC_counter_reg__net3509,
         cu0_counterChain_CounterRC_1_counter_reg__net3515,
         cu0_counterChain_CounterRC_1_counter_reg__net3512,
         cu0_counterChain_CounterRC_1_counter_reg__net3509,
         cu1_counterChain_CounterRC_counter_reg__net3515,
         cu1_counterChain_CounterRC_counter_reg__net3512,
         cu1_counterChain_CounterRC_counter_reg__net3509,
         cu1_counterChain_CounterRC_1_counter_reg__net3518,
         cu1_counterChain_CounterRC_1_counter_reg__net3515,
         cu1_counterChain_CounterRC_1_counter_reg__net3512,
         cu1_counterChain_CounterRC_1_counter_reg__net3509, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345;
  wire   [2:0] cu1_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu1_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu1_RegisterBlock_io_passDataOut_2;
  wire   [6:2] cu1_RegisterBlock_io_passDataOut_3;
  wire   [2:0] cu0_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu0_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu0_RegisterBlock_io_passDataOut_2;
  wire   [7:0] cu0_mem1_mem;
  wire   [7:0] cu1_mem0_mem;
  assign io_status = 1'b0;

  SNPS_CLOCK_GATE_HIGH_SRAM_0_33 cu0_mem1_clk_gate_mem_reg_0_ ( .CLK(clk), 
        .EN(cu0_mem0_N15), .ENCLK(cu0_mem1_net3732), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_32 cu0_mem1_clk_gate_mem_reg_1_ ( .CLK(clk), 
        .EN(cu0_mem0_N16), .ENCLK(cu0_mem1_net3727), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_31 cu0_mem1_clk_gate_mem_reg_2_ ( .CLK(clk), 
        .EN(cu0_mem0_N17), .ENCLK(cu0_mem1_net3722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_30 cu0_mem1_clk_gate_mem_reg_3_ ( .CLK(clk), 
        .EN(cu0_mem0_N18), .ENCLK(cu0_mem1_net3717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_29 cu0_mem1_clk_gate_mem_reg_4_ ( .CLK(clk), 
        .EN(cu0_mem0_N19), .ENCLK(cu0_mem1_net3712), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_28 cu0_mem1_clk_gate_mem_reg_5_ ( .CLK(clk), 
        .EN(cu0_mem0_N20), .ENCLK(cu0_mem1_net3707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_27 cu0_mem1_clk_gate_mem_reg_6_ ( .CLK(clk), 
        .EN(cu0_mem0_N21), .ENCLK(cu0_mem1_net3702), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_26 cu0_mem1_clk_gate_mem_reg_7_ ( .CLK(clk), 
        .EN(cu0_mem0_N22), .ENCLK(cu0_mem1_net3697), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_25 cu0_mem1_clk_gate_mem_reg_8_ ( .CLK(clk), 
        .EN(cu0_mem0_N23), .ENCLK(cu0_mem1_net3692), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_24 cu0_mem1_clk_gate_mem_reg_9_ ( .CLK(clk), 
        .EN(cu0_mem0_N24), .ENCLK(cu0_mem1_net3687), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_23 cu0_mem1_clk_gate_mem_reg_10_ ( .CLK(clk), 
        .EN(cu0_mem0_N25), .ENCLK(cu0_mem1_net3682), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_21 cu0_mem1_clk_gate_mem_reg_12_ ( .CLK(clk), 
        .EN(cu0_mem0_N27), .ENCLK(cu0_mem1_net3672), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_19 cu0_mem1_clk_gate_mem_reg_14_ ( .CLK(clk), 
        .EN(cu0_mem0_N29), .ENCLK(cu0_mem1_net3662), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_18 cu0_mem1_clk_gate_mem_reg_15_ ( .CLK(clk), 
        .EN(cu0_mem0_N30), .ENCLK(cu0_mem1_net3656), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_16 cu1_mem0_clk_gate_mem_reg_0_ ( .CLK(clk), 
        .EN(cu1_mem1_N15), .ENCLK(cu1_mem0_net3732), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_15 cu1_mem0_clk_gate_mem_reg_1_ ( .CLK(clk), 
        .EN(cu1_mem1_N16), .ENCLK(cu1_mem0_net3727), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_14 cu1_mem0_clk_gate_mem_reg_2_ ( .CLK(clk), 
        .EN(cu1_mem1_N17), .ENCLK(cu1_mem0_net3722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_13 cu1_mem0_clk_gate_mem_reg_3_ ( .CLK(clk), 
        .EN(cu1_mem1_N18), .ENCLK(cu1_mem0_net3717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_12 cu1_mem0_clk_gate_mem_reg_4_ ( .CLK(clk), 
        .EN(cu1_mem1_N19), .ENCLK(cu1_mem0_net3712), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_11 cu1_mem0_clk_gate_mem_reg_5_ ( .CLK(clk), 
        .EN(cu1_mem1_N20), .ENCLK(cu1_mem0_net3707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_10 cu1_mem0_clk_gate_mem_reg_6_ ( .CLK(clk), 
        .EN(cu1_mem1_N21), .ENCLK(cu1_mem0_net3702), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_9 cu1_mem0_clk_gate_mem_reg_7_ ( .CLK(clk), .EN(
        cu1_mem1_N22), .ENCLK(cu1_mem0_net3697), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_8 cu1_mem0_clk_gate_mem_reg_8_ ( .CLK(clk), .EN(
        cu1_mem1_N23), .ENCLK(cu1_mem0_net3692), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_7 cu1_mem0_clk_gate_mem_reg_9_ ( .CLK(clk), .EN(
        cu1_mem1_N24), .ENCLK(cu1_mem0_net3687), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_6 cu1_mem0_clk_gate_mem_reg_10_ ( .CLK(clk), 
        .EN(cu1_mem1_N25), .ENCLK(cu1_mem0_net3682), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_4 cu1_mem0_clk_gate_mem_reg_12_ ( .CLK(clk), 
        .EN(cu1_mem1_N27), .ENCLK(cu1_mem0_net3672), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_2 cu1_mem0_clk_gate_mem_reg_14_ ( .CLK(clk), 
        .EN(cu1_mem1_N29), .ENCLK(cu1_mem0_net3662), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_1 cu1_mem0_clk_gate_mem_reg_15_ ( .CLK(clk), 
        .EN(cu1_mem1_N30), .ENCLK(cu1_mem0_net3656), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 cu0_controlBlock_incXbar_clk_gate_config__outSelect_3_reg ( 
        .CLK(clk), .EN(cu0_controlBlock_incXbar_net3599), .ENCLK(
        cu0_controlBlock_incXbar_net3602), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_20 cu0_RegisterBlock_1_FF_1_clk_gate_ff_reg ( 
        .CLK(clk), .EN(cu0_RegisterBlock_1_FF_1_net3491), .ENCLK(
        cu0_RegisterBlock_1_FF_1_net3518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_8 cu1_RegisterBlock_1_FF_1_clk_gate_ff_reg ( 
        .CLK(clk), .EN(cu1_RegisterBlock_1_FF_1_net3491), .ENCLK(
        cu1_RegisterBlock_1_FF_1_net3518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_1 cu1_counterChain_CounterRC_1_counter_reg__clk_gate_ff_reg ( 
        .CLK(clk), .EN(n802), .ENCLK(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .TE(1'b0) );
  DFQD4BWP cu1_controlBlock_config__udcInit_0_reg_1_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_controlBlock_config__udcInit_0_reg_1_ ( .D(n802), .CP(
        cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu1_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu1_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(n802), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(n802), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD1BWP cu1_counterChain_CounterRC_config__stride_reg_0_ ( .D(n802), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_CounterRC_config__stride_0_) );
  DFQD1BWP cu0_config__pipeStage_1_opB_value_reg_0_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net3602), .Q(cu0_T21_0_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3494), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_7_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3494), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_7_) );
  DFQD1BWP controlBox_commandReg_reg ( .D(controlBox_N6), .CP(clk), .Q(
        controlBox_commandReg) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_3_ ( .D(cu0_RegisterBlock_FF_1_net3506), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_3_) );
  DFQD1BWP cu0_mem1_mem_reg_0__0_ ( .D(n1327), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[0]) );
  DFQD1BWP cu0_mem1_mem_reg_0__1_ ( .D(n1326), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[1]) );
  DFQD1BWP cu0_mem1_mem_reg_0__2_ ( .D(n1325), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[2]) );
  DFQD1BWP cu0_mem1_mem_reg_0__3_ ( .D(n1324), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[3]) );
  DFQD1BWP cu0_mem1_mem_reg_0__4_ ( .D(n1323), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[4]) );
  DFQD1BWP cu0_mem1_mem_reg_0__5_ ( .D(n1322), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[5]) );
  DFQD1BWP cu0_mem1_mem_reg_0__6_ ( .D(n1321), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[6]) );
  DFQD1BWP cu0_mem1_mem_reg_0__7_ ( .D(n1320), .CP(cu0_mem1_net3732), .Q(
        cu0_mem1_mem[7]) );
  DFQD1BWP cu1_mem0_mem_reg_0__0_ ( .D(n1335), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[0]) );
  DFQD1BWP cu1_mem0_mem_reg_0__1_ ( .D(n1334), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[1]) );
  DFQD1BWP cu1_mem0_mem_reg_0__2_ ( .D(n1333), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[2]) );
  DFQD1BWP cu1_mem0_mem_reg_0__3_ ( .D(n1332), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[3]) );
  DFQD1BWP cu1_mem0_mem_reg_0__4_ ( .D(n1331), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[4]) );
  DFQD1BWP cu1_mem0_mem_reg_0__5_ ( .D(n1330), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[5]) );
  DFQD1BWP cu1_mem0_mem_reg_0__6_ ( .D(n1329), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[6]) );
  DFQD1BWP cu1_mem0_mem_reg_0__7_ ( .D(n1328), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[7]) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_5_ ( .D(cu0_RegisterBlock_FF_1_net3500), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_6_ ( .D(cu0_RegisterBlock_FF_1_net3497), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_3_ ( .D(cu1_RegisterBlock_FF_1_net3506), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_3_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_5_ ( .D(cu1_RegisterBlock_FF_1_net3500), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_6_ ( .D(cu1_RegisterBlock_FF_1_net3497), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3515), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3512), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3509), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3506), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3503), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3500), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3497), .CP(
        cu0_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3515), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3512), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3509), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3506), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3503), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3500), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_0_ ( .D(cu0_RegisterBlock_FF_1_net3515), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_1_ ( .D(cu0_RegisterBlock_FF_1_net3512), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_2_ ( .D(cu0_RegisterBlock_FF_1_net3509), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_2_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_4_ ( .D(cu0_RegisterBlock_FF_1_net3503), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_2_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3506), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_0_ ( .D(cu1_RegisterBlock_FF_1_net3515), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_0_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_1_ ( .D(cu1_RegisterBlock_FF_1_net3512), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_2_ ( .D(cu1_RegisterBlock_FF_1_net3509), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_4_ ( .D(cu1_RegisterBlock_FF_1_net3503), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(n794) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_0_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3506), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_3_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_4_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_6_) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_3_net3515), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[0]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_3_net3512), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[1]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_3_net3509), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[2]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_3_net3506), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[3]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_3_net3503), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[4]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_3_net3500), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[5]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_3_net3515), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_3_net3512), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[1]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_2_ ( .D(
        cu1_RegisterBlock_FF_3_net3509), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[2]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_3_net3506), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[3]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_3_net3503), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[4]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_3_net3500), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[5]) );
  DFQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .D(
        cu0_counterChain_CounterRC_1_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_1_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_5_ ( .CN(n1336), .D(
        cu1_mem0_mem[5]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[5])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_3_ ( .CN(n1336), .D(
        cu1_mem0_mem[3]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[3])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_0_ ( .CN(n1336), .D(
        cu1_mem0_mem[0]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[0])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_5_ff_reg_6_ ( .CN(n1336), .D(
        cu1_mem0_mem[6]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_3[6])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_5_ff_reg_2_ ( .CN(n1336), .D(
        cu1_mem0_mem[2]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_3[2])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_7_ ( .CN(n1336), .D(
        cu1_mem0_mem[7]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[7])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_4_ ( .CN(n1336), .D(
        cu1_mem0_mem[4]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[4])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_1_ ( .CN(n1336), .D(
        cu1_mem0_mem[1]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[1])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_7_ ( .CN(n1336), .D(
        cu0_mem1_mem[7]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[7])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_6_ ( .CN(n1336), .D(
        cu0_mem1_mem[6]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[6])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_5_ ( .CN(n1336), .D(
        cu0_mem1_mem[5]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[5])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_4_ ( .CN(n1336), .D(
        cu0_mem1_mem[4]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[4])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_3_ ( .CN(n1336), .D(
        cu0_mem1_mem[3]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[3])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_2_ ( .CN(n1336), .D(
        cu0_mem1_mem[2]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[2])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_1_ ( .CN(n1336), .D(
        cu0_mem1_mem[1]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[1])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_0_ ( .CN(n1336), .D(
        cu0_mem1_mem[0]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[0])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_2_ ( .CN(n1336), .D(
        cu1_counterChain_io_data_0_out_2_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[2]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_2_ ( .CN(n1336), .D(
        cu0_counterChain_io_data_0_out_2_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[2]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_1_ ( .CN(n1336), .D(
        cu1_counterChain_io_data_0_out_1_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[1]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_1_ ( .CN(n1336), .D(
        cu0_counterChain_io_data_0_out_1_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[1]) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_0_ ( .CN(n1336), .D(
        cu1_counterChain_io_data_0_out_0_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[0]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_0_ ( .CN(n1336), .D(
        cu0_counterChain_io_data_0_out_0_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[0]) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_0_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_0_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_2_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_2_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_0_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_2_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_1_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_0_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_1_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_2_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_1_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_1_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_6_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_3[6]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_5_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_2_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_3[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_5_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_4_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_3_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_2_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_1_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_0_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_1[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_5_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_4_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_3_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_2_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_1_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_0_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_1[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_7_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_6_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_3[6]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_5_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_4_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_3_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_2_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_3[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_1_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_0_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_7_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_4_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_3_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_1_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_0_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_2_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_0[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_1_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_0[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_0_ ( .CN(n1336), .D(
        cu1_RegisterBlock_io_passDataOut_0[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_7_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_6_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[6]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_5_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_4_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_3_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_2_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_1_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_0_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_7_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_6_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[6]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_5_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_4_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_3_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_2_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_1_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_0_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_2_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_0[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_1_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_0[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_0_ ( .CN(n1336), .D(
        cu0_RegisterBlock_io_passDataOut_0[0]), .CP(clk) );
  DFKCNQD1BWP controlBox_pulser_commandReg_reg ( .CN(n1336), .D(
        controlBox_commandReg), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_0_ ( .CN(n1342), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_0_ ( .CN(n1338), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_7_ ( .CN(n1319), .D(n1337), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_7_ ( .CN(n1319), .D(n1337), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_6_ ( .CN(n1318), .D(n1337), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__0_ ( .CN(1'b1), .D(n1335), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__0_ ( .CN(1'b1), .D(n1327), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_7_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3494), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_7_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3494), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_6_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__1_ ( .CN(1'b1), .D(n1334), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__1_ ( .CN(1'b1), .D(n1326), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_1_ ( .CN(n1343), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_1_ ( .CN(n1339), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__2_ ( .CN(1'b1), .D(n1333), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__2_ ( .CN(1'b1), .D(n1325), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__3_ ( .CN(1'b1), .D(n1332), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__3_ ( .CN(1'b1), .D(n1324), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_2_ ( .CN(n1340), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_2_ ( .CN(n1344), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__4_ ( .CN(1'b1), .D(n1331), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__4_ ( .CN(1'b1), .D(n1323), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__5_ ( .CN(1'b1), .D(n1330), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__5_ ( .CN(1'b1), .D(n1322), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_4_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_4_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_3_ ( .CN(n1341), .D(n1336), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_5_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_5_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_3_ ( .CN(n1336), .D(n1345), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__6_ ( .CN(1'b1), .D(n1329), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__6_ ( .CN(1'b1), .D(n1321), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__7_ ( .CN(1'b1), .D(n1328), .CP(
        cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__7_ ( .CN(1'b1), .D(n1320), .CP(
        cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_7_ ( .CN(n1336), .D(n1328), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_7_ ( .CN(n1336), .D(n1320), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  XOR3D1BWP U972 ( .A1(n783), .A2(n780), .A3(n781), .Z(n786) );
  INR2D1BWP U973 ( .A1(n713), .B1(n685), .ZN(n718) );
  MAOI222D1BWP U974 ( .A(n783), .B(n780), .C(n781), .ZN(n649) );
  CKND1BWP U975 ( .I(n649), .ZN(n711) );
  INR2D1BWP U976 ( .A1(cu1_counterChain_CounterRC_config__stride_0_), .B1(
        reset), .ZN(n834) );
  CKND1BWP U977 ( .I(n795), .ZN(n704) );
  AN2D1BWP U978 ( .A1(n785), .A2(cu0_RegisterBlock_FF_io_data_out_3_), .Z(n797) );
  AO21D1BWP U979 ( .A1(n726), .A2(n727), .B(n731), .Z(n650) );
  OAI211D1BWP U980 ( .A1(n726), .A2(n727), .B(n729), .C(n650), .ZN(n793) );
  CKND2D1BWP U981 ( .A1(cu1_RegisterBlock_1_FF_1_io_data_out_7_), .A2(
        cu0_T21_0_), .ZN(n651) );
  CKXOR2D1BWP U982 ( .A1(n651), .A2(n699), .Z(n1328) );
  CKND2D1BWP U983 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_7_), .A2(
        cu0_T21_0_), .ZN(n652) );
  CKXOR2D1BWP U984 ( .A1(n652), .A2(n678), .Z(n1320) );
  INR2D1BWP U985 ( .A1(n740), .B1(n710), .ZN(n727) );
  IND3D1BWP U986 ( .A1(reset), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n839), .ZN(n842) );
  IND2D1BWP U987 ( .A1(cu0_counterChain_io_data_0_out_2_), .B1(n834), .ZN(n827) );
  AO21D1BWP U988 ( .A1(n664), .A2(n718), .B(n721), .Z(n653) );
  OAI211D1BWP U989 ( .A1(n664), .A2(n718), .B(n729), .C(n653), .ZN(n799) );
  INR2D1BWP U990 ( .A1(n1329), .B1(n802), .ZN(cu1_RegisterBlock_1_FF_1_net3497) );
  INR2D1BWP U991 ( .A1(n1333), .B1(n802), .ZN(cu1_RegisterBlock_1_FF_1_net3509) );
  INR2D1BWP U992 ( .A1(n1321), .B1(n802), .ZN(cu0_RegisterBlock_1_FF_1_net3497) );
  INR2D1BWP U993 ( .A1(n1325), .B1(n802), .ZN(cu0_RegisterBlock_1_FF_1_net3509) );
  IOA21D1BWP U994 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_4_), .B(n690), .ZN(n654) );
  MAOI222D1BWP U995 ( .A(n751), .B(n752), .C(n654), .ZN(n745) );
  XOR3D1BWP U996 ( .A1(n751), .A2(n752), .A3(n654), .Z(n1331) );
  IOA21D1BWP U997 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_4_), .B(n669), .ZN(n655) );
  MAOI222D1BWP U998 ( .A(n753), .B(n754), .C(n655), .ZN(n748) );
  XOR3D1BWP U999 ( .A1(n753), .A2(n754), .A3(n655), .Z(n1323) );
  IND2D1BWP U1000 ( .A1(cu1_counterChain_io_data_0_out_2_), .B1(n834), .ZN(
        n837) );
  ND3D1BWP U1001 ( .A1(cu1_counterChain_CounterRC_config__stride_0_), .A2(n829), .A3(n1336), .ZN(n832) );
  AOI22D1BWP U1002 ( .A1(n777), .A2(n776), .B1(n775), .B2(n774), .ZN(n656) );
  NR2D1BWP U1003 ( .A1(n778), .A2(n656), .ZN(n787) );
  AOI22D1BWP U1004 ( .A1(n783), .A2(n782), .B1(n781), .B2(n780), .ZN(n657) );
  NR2D1BWP U1005 ( .A1(n784), .A2(n657), .ZN(n788) );
  IOA21D1BWP U1006 ( .A1(n785), .A2(n741), .B(n804), .ZN(n1344) );
  IOA21D1BWP U1007 ( .A1(n785), .A2(n714), .B(n803), .ZN(n1340) );
  INR2D1BWP U1008 ( .A1(n1330), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3500) );
  INR2D1BWP U1009 ( .A1(n1331), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3503) );
  INR2D1BWP U1010 ( .A1(n1332), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3506) );
  INR2D1BWP U1011 ( .A1(n1334), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3512) );
  INR2D1BWP U1012 ( .A1(n1335), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3515) );
  INR2D1BWP U1013 ( .A1(n1322), .B1(n802), .ZN(
        cu0_RegisterBlock_1_FF_1_net3500) );
  INR2D1BWP U1014 ( .A1(n1323), .B1(reset), .ZN(
        cu0_RegisterBlock_1_FF_1_net3503) );
  INR2D1BWP U1015 ( .A1(n1324), .B1(reset), .ZN(
        cu0_RegisterBlock_1_FF_1_net3506) );
  INR2D1BWP U1016 ( .A1(n1326), .B1(reset), .ZN(
        cu0_RegisterBlock_1_FF_1_net3512) );
  INR2D1BWP U1017 ( .A1(n1327), .B1(reset), .ZN(
        cu0_RegisterBlock_1_FF_1_net3515) );
  IOA21D1BWP U1018 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_6_), .B(n686), .ZN(n658) );
  MAOI222D1BWP U1019 ( .A(n724), .B(n725), .C(n658), .ZN(n699) );
  XOR3D1BWP U1020 ( .A1(n724), .A2(n725), .A3(n658), .Z(n1329) );
  IOA21D1BWP U1021 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_2_), .B(n694), .ZN(n659) );
  OAI21D1BWP U1022 ( .A1(n785), .A2(n693), .B(n694), .ZN(n660) );
  MAOI222D1BWP U1023 ( .A(n762), .B(n659), .C(n660), .ZN(n758) );
  XOR3D1BWP U1024 ( .A1(n762), .A2(n659), .A3(n660), .Z(n1333) );
  IOA21D1BWP U1025 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_6_), .B(n665), .ZN(n661) );
  MAOI222D1BWP U1026 ( .A(n722), .B(n723), .C(n661), .ZN(n678) );
  XOR3D1BWP U1027 ( .A1(n722), .A2(n723), .A3(n661), .Z(n1321) );
  IOA21D1BWP U1028 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_2_), .B(n673), .ZN(n662) );
  OAI21D1BWP U1029 ( .A1(n785), .A2(n672), .B(n673), .ZN(n663) );
  MAOI222D1BWP U1030 ( .A(n761), .B(n662), .C(n663), .ZN(n755) );
  XOR3D1BWP U1031 ( .A1(n761), .A2(n662), .A3(n663), .Z(n1325) );
  INR2D1BWP U1032 ( .A1(n1328), .B1(n802), .ZN(
        cu1_RegisterBlock_1_FF_1_net3494) );
  INR2D1BWP U1033 ( .A1(n1320), .B1(n802), .ZN(
        cu0_RegisterBlock_1_FF_1_net3494) );
  INVD1BWP U1034 ( .I(cu0_T21_0_), .ZN(n785) );
  AN4D1BWP U1035 ( .A1(n712), .A2(n783), .A3(n780), .A4(n782), .Z(n664) );
  CKND2BWP U1036 ( .I(reset), .ZN(n1336) );
  ND2D1BWP U1487 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_6_), .ZN(
        n665) );
  CKND1BWP U1488 ( .I(n665), .ZN(n723) );
  CKND1BWP U1489 ( .I(cu0_RegisterBlock_io_passDataOut_1[5]), .ZN(n666) );
  ND2D1BWP U1490 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_5_), .ZN(
        n667) );
  OAI21D1BWP U1491 ( .A1(n785), .A2(n666), .B(n667), .ZN(n750) );
  IOA21D1BWP U1492 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_5_), .B(n667), .ZN(n749) );
  CKND1BWP U1493 ( .I(cu0_RegisterBlock_io_passDataOut_1[4]), .ZN(n668) );
  ND2D1BWP U1494 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_4_), .ZN(
        n669) );
  OAI21D1BWP U1495 ( .A1(n785), .A2(n668), .B(n669), .ZN(n754) );
  CKND1BWP U1496 ( .I(cu0_RegisterBlock_io_passDataOut_1[3]), .ZN(n670) );
  ND2D1BWP U1497 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_3_), .ZN(
        n671) );
  OAI21D1BWP U1498 ( .A1(n785), .A2(n670), .B(n671), .ZN(n757) );
  IOA21D1BWP U1499 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_3_), .B(n671), .ZN(n756) );
  CKND1BWP U1500 ( .I(cu0_RegisterBlock_io_passDataOut_1[2]), .ZN(n672) );
  ND2D1BWP U1501 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_2_), .ZN(
        n673) );
  CKND1BWP U1502 ( .I(cu0_RegisterBlock_io_passDataOut_1[1]), .ZN(n674) );
  ND2D1BWP U1503 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_1_), .ZN(
        n675) );
  OAI21D1BWP U1504 ( .A1(n785), .A2(n674), .B(n675), .ZN(n765) );
  IOA21D1BWP U1505 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_1_), .B(n675), .ZN(n764) );
  CKND1BWP U1506 ( .I(cu0_RegisterBlock_io_passDataOut_1[0]), .ZN(n676) );
  ND2D1BWP U1507 ( .A1(n785), .A2(cu0_RegisterBlock_1_FF_io_data_out_0_), .ZN(
        n677) );
  OAI21D1BWP U1508 ( .A1(n785), .A2(n676), .B(n677), .ZN(n771) );
  IOA21D1BWP U1509 ( .A1(cu0_T21_0_), .A2(
        cu0_RegisterBlock_1_FF_1_io_data_out_0_), .B(n677), .ZN(n772) );
  ND2D1BWP U1510 ( .A1(n771), .A2(n772), .ZN(n763) );
  CKND2D1BWP U1511 ( .A1(n785), .A2(cu0_RegisterBlock_FF_io_data_out_2_), .ZN(
        n679) );
  IOA21D1BWP U1512 ( .A1(cu0_T21_0_), .A2(cu0_counterChain_io_data_1_out_2_), 
        .B(n679), .ZN(n712) );
  CKND1BWP U1513 ( .I(n712), .ZN(n685) );
  IOA21D1BWP U1514 ( .A1(cu0_T21_0_), .A2(cu0_counterChain_io_data_0_out_2_), 
        .B(n679), .ZN(n713) );
  INVD1BWP U1515 ( .I(cu0_counterChain_io_data_1_out_1_), .ZN(n831) );
  ND2D1BWP U1516 ( .A1(n785), .A2(cu0_RegisterBlock_FF_io_data_out_1_), .ZN(
        n680) );
  OAI21D1BWP U1517 ( .A1(n785), .A2(n831), .B(n680), .ZN(n783) );
  AN2XD1BWP U1518 ( .A1(n783), .A2(n713), .Z(n702) );
  CKND1BWP U1519 ( .I(cu0_counterChain_io_data_1_out_0_), .ZN(n830) );
  CKND2D1BWP U1520 ( .A1(n785), .A2(cu0_RegisterBlock_FF_io_data_out_0_), .ZN(
        n681) );
  OAI21D1BWP U1521 ( .A1(n830), .A2(n785), .B(n681), .ZN(n781) );
  INVD1BWP U1522 ( .I(cu0_counterChain_io_data_0_out_1_), .ZN(n826) );
  OAI21D1BWP U1523 ( .A1(n785), .A2(n826), .B(n680), .ZN(n780) );
  CKND1BWP U1524 ( .I(cu0_counterChain_io_data_0_out_0_), .ZN(n825) );
  OAI21D1BWP U1525 ( .A1(n825), .A2(n785), .B(n681), .ZN(n782) );
  AN4D1BWP U1526 ( .A1(n783), .A2(n781), .A3(n780), .A4(n782), .Z(n784) );
  CKND1BWP U1527 ( .I(n782), .ZN(n683) );
  CKND2D1BWP U1528 ( .A1(n783), .A2(n780), .ZN(n682) );
  OAI32D1BWP U1529 ( .A1(n664), .A2(n685), .A3(n683), .B1(n682), .B2(n664), 
        .ZN(n716) );
  AN2XD1BWP U1530 ( .A1(n781), .A2(n713), .Z(n715) );
  CKND1BWP U1531 ( .I(n780), .ZN(n684) );
  AOI211D1BWP U1532 ( .A1(n783), .A2(n782), .B(n685), .C(n684), .ZN(n700) );
  NR2D1BWP U1533 ( .A1(n785), .A2(reset), .ZN(n729) );
  CKND1BWP U1534 ( .I(n799), .ZN(cu0_RegisterBlock_FF_3_net3500) );
  ND2D1BWP U1535 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_6_), .ZN(
        n686) );
  CKND1BWP U1536 ( .I(n686), .ZN(n725) );
  CKND1BWP U1537 ( .I(cu1_RegisterBlock_io_passDataOut_1[5]), .ZN(n687) );
  ND2D1BWP U1538 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_5_), .ZN(
        n688) );
  OAI21D1BWP U1539 ( .A1(n785), .A2(n687), .B(n688), .ZN(n747) );
  IOA21D1BWP U1540 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_5_), .B(n688), .ZN(n746) );
  CKND1BWP U1541 ( .I(cu1_RegisterBlock_io_passDataOut_1[4]), .ZN(n689) );
  ND2D1BWP U1542 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_4_), .ZN(
        n690) );
  OAI21D1BWP U1543 ( .A1(n785), .A2(n689), .B(n690), .ZN(n752) );
  CKND1BWP U1544 ( .I(cu1_RegisterBlock_io_passDataOut_1[3]), .ZN(n691) );
  ND2D1BWP U1545 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_3_), .ZN(
        n692) );
  OAI21D1BWP U1546 ( .A1(n785), .A2(n691), .B(n692), .ZN(n760) );
  IOA21D1BWP U1547 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_3_), .B(n692), .ZN(n759) );
  CKND1BWP U1548 ( .I(cu1_RegisterBlock_io_passDataOut_1[2]), .ZN(n693) );
  ND2D1BWP U1549 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_2_), .ZN(
        n694) );
  CKND1BWP U1550 ( .I(cu1_RegisterBlock_io_passDataOut_1[1]), .ZN(n695) );
  ND2D1BWP U1551 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_1_), .ZN(
        n696) );
  OAI21D1BWP U1552 ( .A1(n785), .A2(n695), .B(n696), .ZN(n768) );
  IOA21D1BWP U1553 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_1_), .B(n696), .ZN(n767) );
  CKND1BWP U1554 ( .I(cu1_RegisterBlock_io_passDataOut_1[0]), .ZN(n697) );
  ND2D1BWP U1555 ( .A1(n785), .A2(cu1_RegisterBlock_1_FF_io_data_out_0_), .ZN(
        n698) );
  OAI21D1BWP U1556 ( .A1(n785), .A2(n697), .B(n698), .ZN(n769) );
  IOA21D1BWP U1557 ( .A1(cu0_T21_0_), .A2(
        cu1_RegisterBlock_1_FF_1_io_data_out_0_), .B(n698), .ZN(n770) );
  ND2D1BWP U1558 ( .A1(n769), .A2(n770), .ZN(n766) );
  FA1D1BWP U1559 ( .A(n702), .B(n701), .CI(n700), .CO(n721), .S(n703) );
  CKND2D1BWP U1560 ( .A1(cu0_T21_0_), .A2(n703), .ZN(n792) );
  IOA21D1BWP U1561 ( .A1(n704), .A2(n785), .B(n792), .ZN(n1341) );
  CKND2D1BWP U1562 ( .A1(n785), .A2(cu1_RegisterBlock_FF_io_data_out_2_), .ZN(
        n705) );
  IOA21D1BWP U1563 ( .A1(cu0_T21_0_), .A2(cu1_counterChain_io_data_1_out_2_), 
        .B(n705), .ZN(n739) );
  CKND1BWP U1564 ( .I(n739), .ZN(n710) );
  IOA21D1BWP U1565 ( .A1(cu0_T21_0_), .A2(cu1_counterChain_io_data_0_out_2_), 
        .B(n705), .ZN(n740) );
  INVD1BWP U1566 ( .I(cu1_counterChain_io_data_1_out_1_), .ZN(n841) );
  ND2D1BWP U1567 ( .A1(n785), .A2(cu1_RegisterBlock_FF_io_data_out_1_), .ZN(
        n706) );
  OAI21D1BWP U1568 ( .A1(n785), .A2(n841), .B(n706), .ZN(n777) );
  AN2XD1BWP U1569 ( .A1(n777), .A2(n740), .Z(n735) );
  CKND1BWP U1570 ( .I(cu1_counterChain_io_data_1_out_0_), .ZN(n840) );
  CKND2D1BWP U1571 ( .A1(n785), .A2(cu1_RegisterBlock_FF_io_data_out_0_), .ZN(
        n707) );
  OAI21D1BWP U1572 ( .A1(n840), .A2(n785), .B(n707), .ZN(n775) );
  INVD1BWP U1573 ( .I(cu1_counterChain_io_data_0_out_1_), .ZN(n836) );
  OAI21D1BWP U1574 ( .A1(n785), .A2(n836), .B(n706), .ZN(n774) );
  CKND1BWP U1575 ( .I(cu1_counterChain_io_data_0_out_0_), .ZN(n835) );
  OAI21D1BWP U1576 ( .A1(n835), .A2(n785), .B(n707), .ZN(n776) );
  AN4D1BWP U1577 ( .A1(n777), .A2(n775), .A3(n774), .A4(n776), .Z(n778) );
  AN4D1BWP U1578 ( .A1(n739), .A2(n777), .A3(n774), .A4(n776), .Z(n726) );
  CKND1BWP U1579 ( .I(n776), .ZN(n773) );
  CKND2D1BWP U1580 ( .A1(n777), .A2(n774), .ZN(n708) );
  OAI32D1BWP U1581 ( .A1(n726), .A2(n710), .A3(n773), .B1(n708), .B2(n726), 
        .ZN(n743) );
  AN2XD1BWP U1582 ( .A1(n775), .A2(n740), .Z(n742) );
  CKND1BWP U1583 ( .I(n774), .ZN(n709) );
  AOI211D1BWP U1584 ( .A1(n777), .A2(n776), .B(n710), .C(n709), .ZN(n733) );
  CKND1BWP U1585 ( .I(n793), .ZN(cu1_RegisterBlock_FF_3_net3500) );
  FICOND1BWP U1586 ( .A(n713), .B(n712), .CI(n711), .CON(n795), .S(n714) );
  FA1D1BWP U1587 ( .A(n784), .B(n716), .CI(n715), .CO(n701), .S(n717) );
  CKND2D1BWP U1588 ( .A1(cu0_T21_0_), .A2(n717), .ZN(n803) );
  MAOI22D1BWP U1589 ( .A1(n718), .A2(n664), .B1(n664), .B2(n718), .ZN(n720) );
  ND2D1BWP U1590 ( .A1(n721), .A2(n720), .ZN(n719) );
  OAI211D1BWP U1591 ( .A1(n721), .A2(n720), .B(n729), .C(n719), .ZN(n796) );
  CKND1BWP U1592 ( .I(n796), .ZN(cu0_RegisterBlock_FF_3_net3503) );
  MAOI22D1BWP U1593 ( .A1(n727), .A2(n726), .B1(n726), .B2(n727), .ZN(n730) );
  ND2D1BWP U1594 ( .A1(n731), .A2(n730), .ZN(n728) );
  OAI211D1BWP U1595 ( .A1(n731), .A2(n730), .B(n729), .C(n728), .ZN(n791) );
  CKND1BWP U1596 ( .I(n791), .ZN(cu1_RegisterBlock_FF_3_net3503) );
  CKND2D1BWP U1597 ( .A1(n732), .A2(n785), .ZN(n737) );
  FA1D1BWP U1598 ( .A(n735), .B(n734), .CI(n733), .CO(n731), .S(n736) );
  CKND2D1BWP U1599 ( .A1(cu0_T21_0_), .A2(n736), .ZN(n789) );
  ND2D1BWP U1600 ( .A1(n737), .A2(n789), .ZN(n1345) );
  FICOND1BWP U1601 ( .A(n740), .B(n739), .CI(n738), .CON(n790), .S(n741) );
  FA1D1BWP U1602 ( .A(n778), .B(n743), .CI(n742), .CO(n734), .S(n744) );
  CKND2D1BWP U1603 ( .A1(cu0_T21_0_), .A2(n744), .ZN(n804) );
  FICIND1BWP U1604 ( .CIN(n745), .B(n746), .A(n747), .CO(n724), .S(n1330) );
  FICIND1BWP U1605 ( .CIN(n748), .B(n749), .A(n750), .CO(n722), .S(n1322) );
  FICIND1BWP U1606 ( .CIN(n755), .B(n756), .A(n757), .CO(n753), .S(n1324) );
  FICIND1BWP U1607 ( .CIN(n758), .B(n759), .A(n760), .CO(n751), .S(n1332) );
  NR2D1BWP U1608 ( .A1(cu0_T21_0_), .A2(reset), .ZN(n800) );
  CKND1BWP U1609 ( .I(cu0_RegisterBlock_FF_io_data_out_4_), .ZN(n798) );
  AN2XD1BWP U1610 ( .A1(n800), .A2(cu0_RegisterBlock_FF_io_data_out_6_), .Z(
        cu0_RegisterBlock_FF_1_net3494) );
  FICIND1BWP U1611 ( .CIN(n763), .B(n764), .A(n765), .CO(n761), .S(n1326) );
  FICIND1BWP U1612 ( .CIN(n766), .B(n767), .A(n768), .CO(n762), .S(n1334) );
  XOR2D1BWP U1613 ( .A1(n770), .A2(n769), .Z(n1335) );
  AN2XD1BWP U1614 ( .A1(n800), .A2(cu0_RegisterBlock_FF_io_data_out_5_), .Z(
        cu0_RegisterBlock_FF_1_net3497) );
  XOR2D1BWP U1615 ( .A1(n772), .A2(n771), .Z(n1327) );
  NR2D1BWP U1616 ( .A1(n802), .A2(cu0_T21_0_), .ZN(n1337) );
  CKAN2D1BWP U1617 ( .A1(n785), .A2(cu1_RegisterBlock_FF_io_data_out_5_), .Z(
        n1318) );
  AN2XD1BWP U1618 ( .A1(n1337), .A2(n1318), .Z(cu1_RegisterBlock_FF_1_net3497)
         );
  CKND1BWP U1619 ( .I(n800), .ZN(cu0_RegisterBlock_1_FF_1_net3491) );
  CKND1BWP U1620 ( .I(n1337), .ZN(cu1_RegisterBlock_1_FF_1_net3491) );
  ND3D1BWP U1621 ( .A1(cu0_counterChain_io_data_0_out_0_), .A2(
        cu0_counterChain_io_data_1_out_0_), .A3(cu0_T21_0_), .ZN(n845) );
  CKND1BWP U1622 ( .I(n845), .ZN(n1338) );
  ND3D1BWP U1623 ( .A1(cu1_counterChain_io_data_1_out_0_), .A2(
        cu1_counterChain_io_data_0_out_0_), .A3(cu0_T21_0_), .ZN(n857) );
  CKND1BWP U1624 ( .I(n857), .ZN(n1342) );
  OR2XD1BWP U1625 ( .A1(io_config_enable), .A2(n802), .Z(
        cu0_controlBlock_incXbar_net3599) );
  CKAN2D1BWP U1626 ( .A1(n785), .A2(cu1_RegisterBlock_FF_io_data_out_6_), .Z(
        n1319) );
  FICIND1BWP U1627 ( .CIN(n773), .B(n777), .A(n774), .CO(n738), .S(n779) );
  AO21D1BWP U1628 ( .A1(n779), .A2(n785), .B(n787), .Z(n1343) );
  AO21D1BWP U1629 ( .A1(n786), .A2(n785), .B(n788), .Z(n1339) );
  NR2D1BWP U1630 ( .A1(reset), .A2(n857), .ZN(cu1_RegisterBlock_FF_1_net3515)
         );
  NR2D1BWP U1631 ( .A1(n802), .A2(n845), .ZN(cu0_RegisterBlock_FF_1_net3515)
         );
  MOAI22D1BWP U1632 ( .A1(n841), .A2(cu1_RegisterBlock_1_FF_1_net3491), .B1(
        n1336), .B2(n787), .ZN(cu1_RegisterBlock_FF_3_net3512) );
  INVD1BWP U1633 ( .I(n1336), .ZN(n802) );
  MOAI22D1BWP U1634 ( .A1(n831), .A2(cu0_RegisterBlock_1_FF_1_net3491), .B1(
        n1336), .B2(n788), .ZN(cu0_RegisterBlock_FF_3_net3512) );
  INVD1BWP U1635 ( .I(n1343), .ZN(n856) );
  NR2D1BWP U1636 ( .A1(reset), .A2(n856), .ZN(cu1_RegisterBlock_FF_1_net3512)
         );
  INVD1BWP U1637 ( .I(n1339), .ZN(n844) );
  NR2D1BWP U1638 ( .A1(reset), .A2(n844), .ZN(cu0_RegisterBlock_FF_1_net3512)
         );
  CKND1BWP U1639 ( .I(n1344), .ZN(n861) );
  NR2D1BWP U1640 ( .A1(reset), .A2(n861), .ZN(cu1_RegisterBlock_FF_1_net3509)
         );
  NR2D1BWP U1641 ( .A1(reset), .A2(n789), .ZN(cu1_RegisterBlock_FF_3_net3506)
         );
  CKND1BWP U1642 ( .I(n1340), .ZN(n849) );
  NR2D1BWP U1643 ( .A1(n802), .A2(n849), .ZN(cu0_RegisterBlock_FF_1_net3509)
         );
  FICIND1BWP U1644 ( .CIN(n790), .B(cu1_RegisterBlock_FF_io_data_out_3_), .A(
        cu1_RegisterBlock_FF_io_data_out_3_), .S(n732) );
  IOA21D1BWP U1645 ( .A1(cu1_RegisterBlock_FF_io_data_out_3_), .A2(n1337), .B(
        n791), .ZN(cu1_RegisterBlock_FF_1_net3503) );
  NR2D1BWP U1646 ( .A1(n802), .A2(n792), .ZN(cu0_RegisterBlock_FF_3_net3506)
         );
  IOA21D1BWP U1647 ( .A1(n794), .A2(n1337), .B(n793), .ZN(
        cu1_RegisterBlock_FF_1_net3500) );
  CKND1BWP U1648 ( .I(n1345), .ZN(n859) );
  NR2D1BWP U1649 ( .A1(n859), .A2(n802), .ZN(cu1_RegisterBlock_FF_1_net3506)
         );
  IOA21D1BWP U1650 ( .A1(n797), .A2(n800), .B(n796), .ZN(
        cu0_RegisterBlock_FF_1_net3503) );
  FICIND1BWP U1651 ( .CIN(n798), .B(cu0_RegisterBlock_FF_io_data_out_5_), .A(
        cu0_RegisterBlock_FF_io_data_out_5_), .S(n801) );
  IOA21D1BWP U1652 ( .A1(n801), .A2(n800), .B(n799), .ZN(
        cu0_RegisterBlock_FF_1_net3500) );
  CKND1BWP U1653 ( .I(n1341), .ZN(n847) );
  NR2D1BWP U1654 ( .A1(reset), .A2(n847), .ZN(cu0_RegisterBlock_FF_1_net3506)
         );
  AOI211D1BWP U1656 ( .A1(cu0_T21_0_), .A2(n825), .B(n802), .C(n830), .ZN(
        cu0_RegisterBlock_FF_3_net3515) );
  CKND1BWP U1657 ( .I(cu0_counterChain_io_data_1_out_2_), .ZN(n829) );
  OAI22D1BWP U1658 ( .A1(n802), .A2(n803), .B1(n829), .B2(
        cu0_RegisterBlock_1_FF_1_net3491), .ZN(cu0_RegisterBlock_FF_3_net3509)
         );
  AOI211D1BWP U1659 ( .A1(cu0_T21_0_), .A2(n835), .B(reset), .C(n840), .ZN(
        cu1_RegisterBlock_FF_3_net3515) );
  CKND1BWP U1660 ( .I(cu1_counterChain_io_data_1_out_2_), .ZN(n839) );
  OAI22D1BWP U1661 ( .A1(reset), .A2(n804), .B1(n839), .B2(
        cu1_RegisterBlock_1_FF_1_net3491), .ZN(cu1_RegisterBlock_FF_3_net3509)
         );
  NR2D1BWP U1662 ( .A1(reset), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3581) );
  INR2D1BWP U1663 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__net3581), .B1(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n805) );
  AO31D1BWP U1664 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), 
        .A2(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n1336), .B(
        n805), .Z(cu1_controlBlock_UpDownCtr_1_reg__net3578) );
  NR2D1BWP U1665 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n807) );
  CKND1BWP U1666 ( .I(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n806) );
  ND2D1BWP U1667 ( .A1(n805), .A2(n806), .ZN(n809) );
  OAI31D1BWP U1668 ( .A1(reset), .A2(n807), .A3(n806), .B(n809), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3575) );
  OAI31D1BWP U1669 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n808) );
  OAI22D1BWP U1670 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n809), .B1(n802), .B2(n808), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3572) );
  NR2D1BWP U1671 ( .A1(n802), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3581) );
  INR2D1BWP U1672 ( .A1(cu0_controlBlock_UpDownCtr_reg__net3581), .B1(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n810) );
  AO31D1BWP U1673 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n1336), .B(n810), 
        .Z(cu0_controlBlock_UpDownCtr_reg__net3578) );
  NR2D1BWP U1674 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n812) );
  CKND1BWP U1675 ( .I(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(
        n811) );
  ND2D1BWP U1676 ( .A1(n810), .A2(n811), .ZN(n814) );
  OAI31D1BWP U1677 ( .A1(reset), .A2(n812), .A3(n811), .B(n814), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3575) );
  OAI31D1BWP U1678 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n813) );
  OAI22D1BWP U1679 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n814), .B1(reset), .B2(n813), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3572) );
  NR2D1BWP U1680 ( .A1(reset), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3581) );
  INR2D1BWP U1681 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__net3581), .B1(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n815) );
  AO31D1BWP U1682 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), 
        .A2(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n1336), .B(
        n815), .Z(cu0_controlBlock_UpDownCtr_1_reg__net3578) );
  NR2D1BWP U1683 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n817) );
  CKND1BWP U1684 ( .I(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n816) );
  ND2D1BWP U1685 ( .A1(n815), .A2(n816), .ZN(n819) );
  OAI31D1BWP U1686 ( .A1(reset), .A2(n817), .A3(n816), .B(n819), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3575) );
  OAI31D1BWP U1687 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n818) );
  OAI22D1BWP U1688 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n819), .B1(n802), .B2(n818), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3572) );
  NR2D1BWP U1689 ( .A1(n802), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3581) );
  INR2D1BWP U1690 ( .A1(cu1_controlBlock_UpDownCtr_reg__net3581), .B1(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n820) );
  AO31D1BWP U1691 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n1336), .B(n820), 
        .Z(cu1_controlBlock_UpDownCtr_reg__net3578) );
  NR2D1BWP U1692 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n822) );
  CKND1BWP U1693 ( .I(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(
        n821) );
  ND2D1BWP U1694 ( .A1(n820), .A2(n821), .ZN(n824) );
  OAI31D1BWP U1695 ( .A1(reset), .A2(n822), .A3(n821), .B(n824), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3575) );
  OAI31D1BWP U1696 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n823) );
  OAI22D1BWP U1697 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n824), .B1(reset), .B2(n823), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3572) );
  NR2D1BWP U1698 ( .A1(n827), .A2(cu0_counterChain_io_data_0_out_0_), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net3515) );
  AOI221D1BWP U1699 ( .A1(cu0_counterChain_io_data_0_out_1_), .A2(
        cu0_counterChain_io_data_0_out_0_), .B1(n826), .B2(n825), .C(n827), 
        .ZN(cu0_counterChain_CounterRC_counter_reg__net3512) );
  CKND2D1BWP U1700 ( .A1(cu0_counterChain_io_data_0_out_1_), .A2(
        cu0_counterChain_io_data_0_out_0_), .ZN(n828) );
  NR2D1BWP U1701 ( .A1(n828), .A2(n827), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net3509) );
  NR2D1BWP U1702 ( .A1(n832), .A2(cu0_counterChain_io_data_1_out_0_), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net3515) );
  AOI221D1BWP U1703 ( .A1(cu0_counterChain_io_data_1_out_1_), .A2(
        cu0_counterChain_io_data_1_out_0_), .B1(n831), .B2(n830), .C(n832), 
        .ZN(cu0_counterChain_CounterRC_1_counter_reg__net3512) );
  CKND2D1BWP U1704 ( .A1(cu0_counterChain_io_data_1_out_1_), .A2(
        cu0_counterChain_io_data_1_out_0_), .ZN(n833) );
  NR2D1BWP U1705 ( .A1(n833), .A2(n832), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net3509) );
  NR2D1BWP U1706 ( .A1(n837), .A2(cu1_counterChain_io_data_0_out_0_), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net3515) );
  AOI221D1BWP U1707 ( .A1(cu1_counterChain_io_data_0_out_1_), .A2(
        cu1_counterChain_io_data_0_out_0_), .B1(n836), .B2(n835), .C(n837), 
        .ZN(cu1_counterChain_CounterRC_counter_reg__net3512) );
  CKND2D1BWP U1708 ( .A1(cu1_counterChain_io_data_0_out_1_), .A2(
        cu1_counterChain_io_data_0_out_0_), .ZN(n838) );
  NR2D1BWP U1709 ( .A1(n838), .A2(n837), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net3509) );
  NR2D1BWP U1710 ( .A1(n842), .A2(cu1_counterChain_io_data_1_out_0_), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net3515) );
  AOI221D1BWP U1711 ( .A1(cu1_counterChain_io_data_1_out_1_), .A2(
        cu1_counterChain_io_data_1_out_0_), .B1(n841), .B2(n840), .C(n842), 
        .ZN(cu1_counterChain_CounterRC_1_counter_reg__net3512) );
  CKND2D1BWP U1712 ( .A1(cu1_counterChain_io_data_1_out_1_), .A2(
        cu1_counterChain_io_data_1_out_0_), .ZN(n843) );
  NR2D1BWP U1713 ( .A1(n843), .A2(n842), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net3509) );
  ND2D1BWP U1714 ( .A1(n847), .A2(n849), .ZN(n846) );
  ND2D1BWP U1715 ( .A1(n844), .A2(n845), .ZN(n852) );
  NR2D1BWP U1716 ( .A1(n846), .A2(n852), .ZN(cu0_mem0_N15) );
  ND2D1BWP U1717 ( .A1(n844), .A2(n1338), .ZN(n850) );
  NR2D1BWP U1718 ( .A1(n850), .A2(n846), .ZN(cu0_mem0_N16) );
  ND2D1BWP U1719 ( .A1(n1339), .A2(n845), .ZN(n853) );
  NR2D1BWP U1720 ( .A1(n853), .A2(n846), .ZN(cu0_mem0_N17) );
  ND2D1BWP U1721 ( .A1(n1339), .A2(n1338), .ZN(n854) );
  NR2D1BWP U1722 ( .A1(n854), .A2(n846), .ZN(cu0_mem0_N18) );
  ND2D1BWP U1723 ( .A1(n847), .A2(n1340), .ZN(n848) );
  NR2D1BWP U1724 ( .A1(n848), .A2(n852), .ZN(cu0_mem0_N19) );
  NR2D1BWP U1725 ( .A1(n848), .A2(n850), .ZN(cu0_mem0_N20) );
  NR2D1BWP U1726 ( .A1(n848), .A2(n853), .ZN(cu0_mem0_N21) );
  NR2D1BWP U1727 ( .A1(n848), .A2(n854), .ZN(cu0_mem0_N22) );
  CKND2D1BWP U1728 ( .A1(n1341), .A2(n849), .ZN(n851) );
  NR2D1BWP U1729 ( .A1(n851), .A2(n852), .ZN(cu0_mem0_N23) );
  NR2D1BWP U1730 ( .A1(n851), .A2(n850), .ZN(cu0_mem0_N24) );
  NR2D1BWP U1731 ( .A1(n851), .A2(n853), .ZN(cu0_mem0_N25) );
  CKND2D1BWP U1732 ( .A1(n1341), .A2(n1340), .ZN(n855) );
  NR2D1BWP U1733 ( .A1(n855), .A2(n852), .ZN(cu0_mem0_N27) );
  NR2D1BWP U1734 ( .A1(n855), .A2(n853), .ZN(cu0_mem0_N29) );
  NR2D1BWP U1735 ( .A1(n855), .A2(n854), .ZN(cu0_mem0_N30) );
  ND2D1BWP U1736 ( .A1(n859), .A2(n861), .ZN(n858) );
  ND2D1BWP U1737 ( .A1(n856), .A2(n857), .ZN(n864) );
  NR2D1BWP U1738 ( .A1(n858), .A2(n864), .ZN(cu1_mem1_N15) );
  ND2D1BWP U1739 ( .A1(n856), .A2(n1342), .ZN(n862) );
  NR2D1BWP U1740 ( .A1(n862), .A2(n858), .ZN(cu1_mem1_N16) );
  ND2D1BWP U1741 ( .A1(n1343), .A2(n857), .ZN(n865) );
  NR2D1BWP U1742 ( .A1(n865), .A2(n858), .ZN(cu1_mem1_N17) );
  ND2D1BWP U1743 ( .A1(n1343), .A2(n1342), .ZN(n866) );
  NR2D1BWP U1744 ( .A1(n866), .A2(n858), .ZN(cu1_mem1_N18) );
  ND2D1BWP U1745 ( .A1(n859), .A2(n1344), .ZN(n860) );
  NR2D1BWP U1746 ( .A1(n860), .A2(n864), .ZN(cu1_mem1_N19) );
  NR2D1BWP U1747 ( .A1(n860), .A2(n862), .ZN(cu1_mem1_N20) );
  NR2D1BWP U1748 ( .A1(n860), .A2(n865), .ZN(cu1_mem1_N21) );
  NR2D1BWP U1749 ( .A1(n860), .A2(n866), .ZN(cu1_mem1_N22) );
  CKND2D1BWP U1750 ( .A1(n1345), .A2(n861), .ZN(n863) );
  NR2D1BWP U1751 ( .A1(n863), .A2(n864), .ZN(cu1_mem1_N23) );
  NR2D1BWP U1752 ( .A1(n863), .A2(n862), .ZN(cu1_mem1_N24) );
  NR2D1BWP U1753 ( .A1(n863), .A2(n865), .ZN(cu1_mem1_N25) );
  CKND2D1BWP U1754 ( .A1(n1345), .A2(n1344), .ZN(n867) );
  NR2D1BWP U1755 ( .A1(n867), .A2(n864), .ZN(cu1_mem1_N27) );
  NR2D1BWP U1756 ( .A1(n867), .A2(n865), .ZN(cu1_mem1_N29) );
  NR2D1BWP U1757 ( .A1(n867), .A2(n866), .ZN(cu1_mem1_N30) );
  INR2D1BWP U1758 ( .A1(io_command), .B1(n802), .ZN(controlBox_N6) );
endmodule

