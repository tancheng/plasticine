
module SNPS_CLOCK_GATE_HIGH_FF_1_4_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FF_1_4_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_SRAM_0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module Plasticine ( clk, reset, io_config_enable, io_command, io_status );
  input clk, reset, io_config_enable, io_command;
  output io_status;
  wire   controlBox_N6, controlBox_commandReg,
         cu1_RegisterBlock_io_passDataOut_3_6_,
         cu1_counterChain_io_data_0_out_0_, cu1_counterChain_io_data_0_out_1_,
         cu1_counterChain_io_data_0_out_2_, cu1_counterChain_io_data_1_out_0_,
         cu1_counterChain_io_data_1_out_1_, cu1_counterChain_io_data_1_out_2_,
         cu0_counterChain_io_data_0_out_0_, cu0_counterChain_io_data_0_out_1_,
         cu0_counterChain_io_data_0_out_2_, cu0_counterChain_io_data_1_out_0_,
         cu0_counterChain_io_data_1_out_1_, cu0_counterChain_io_data_1_out_2_,
         cu1_mem1_N30, cu1_mem1_N29, cu1_mem1_N27, cu1_mem1_N25, cu1_mem1_N24,
         cu1_mem1_N23, cu1_mem1_N22, cu1_mem1_N21, cu1_mem1_N20, cu1_mem1_N19,
         cu1_mem1_N18, cu1_mem1_N17, cu1_mem1_N16, cu1_mem1_N15,
         cu1_mem1_mem_0__6_, cu1_RegisterBlock_1_FF_1_io_data_out_0_,
         cu1_RegisterBlock_1_FF_1_io_data_out_1_,
         cu1_RegisterBlock_1_FF_1_io_data_out_2_,
         cu1_RegisterBlock_1_FF_1_io_data_out_3_,
         cu1_RegisterBlock_1_FF_1_io_data_out_4_,
         cu1_RegisterBlock_1_FF_1_io_data_out_5_,
         cu1_RegisterBlock_1_FF_1_io_data_out_6_,
         cu1_RegisterBlock_1_FF_1_io_data_out_7_,
         cu1_RegisterBlock_1_FF_io_data_out_0_,
         cu1_RegisterBlock_1_FF_io_data_out_1_,
         cu1_RegisterBlock_1_FF_io_data_out_2_,
         cu1_RegisterBlock_1_FF_io_data_out_3_,
         cu1_RegisterBlock_1_FF_io_data_out_4_,
         cu1_RegisterBlock_1_FF_io_data_out_5_,
         cu1_RegisterBlock_1_FF_io_data_out_6_,
         cu1_RegisterBlock_FF_io_data_out_0_,
         cu1_RegisterBlock_FF_io_data_out_1_,
         cu1_RegisterBlock_FF_io_data_out_2_,
         cu1_RegisterBlock_FF_io_data_out_3_,
         cu1_RegisterBlock_FF_io_data_out_4_,
         cu1_RegisterBlock_FF_io_data_out_5_,
         cu1_RegisterBlock_FF_io_data_out_6_, cu0_mem0_N30, cu0_mem0_N29,
         cu0_mem0_N27, cu0_mem0_N25, cu0_mem0_N24, cu0_mem0_N23, cu0_mem0_N22,
         cu0_mem0_N21, cu0_mem0_N20, cu0_mem0_N19, cu0_mem0_N18, cu0_mem0_N17,
         cu0_mem0_N16, cu0_mem0_N15, cu0_mem1_net3732, cu0_mem1_net3727,
         cu0_mem1_net3722, cu0_mem1_net3717, cu0_mem1_net3712,
         cu0_mem1_net3707, cu0_mem1_net3702, cu0_mem1_net3697,
         cu0_mem1_net3692, cu0_mem1_net3687, cu0_mem1_net3682,
         cu0_mem1_net3672, cu0_mem1_net3662, cu0_mem1_net3656,
         cu0_RegisterBlock_FF_io_data_out_0_,
         cu0_RegisterBlock_FF_io_data_out_1_,
         cu0_RegisterBlock_FF_io_data_out_2_,
         cu0_RegisterBlock_FF_io_data_out_3_,
         cu0_RegisterBlock_FF_io_data_out_4_,
         cu0_RegisterBlock_FF_io_data_out_5_,
         cu0_RegisterBlock_FF_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_0_,
         cu0_RegisterBlock_1_FF_1_io_data_out_1_,
         cu0_RegisterBlock_1_FF_1_io_data_out_2_,
         cu0_RegisterBlock_1_FF_1_io_data_out_3_,
         cu0_RegisterBlock_1_FF_1_io_data_out_4_,
         cu0_RegisterBlock_1_FF_1_io_data_out_5_,
         cu0_RegisterBlock_1_FF_1_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_7_,
         cu0_RegisterBlock_1_FF_io_data_out_0_,
         cu0_RegisterBlock_1_FF_io_data_out_1_,
         cu0_RegisterBlock_1_FF_io_data_out_2_,
         cu0_RegisterBlock_1_FF_io_data_out_3_,
         cu0_RegisterBlock_1_FF_io_data_out_4_,
         cu0_RegisterBlock_1_FF_io_data_out_5_,
         cu0_RegisterBlock_1_FF_io_data_out_6_, cu1_mem0_net3732,
         cu1_mem0_net3727, cu1_mem0_net3722, cu1_mem0_net3717,
         cu1_mem0_net3712, cu1_mem0_net3707, cu1_mem0_net3702,
         cu1_mem0_net3697, cu1_mem0_net3692, cu1_mem0_net3687,
         cu1_mem0_net3682, cu1_mem0_net3672, cu1_mem0_net3662,
         cu1_mem0_net3656, cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_incXbar_net3602, cu0_controlBlock_incXbar_net3599,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu0_RegisterBlock_FF_1_net3506, cu0_RegisterBlock_FF_1_net3503,
         cu0_RegisterBlock_FF_1_net3500, cu0_RegisterBlock_FF_1_net3497,
         cu0_RegisterBlock_FF_3_net3515, cu0_RegisterBlock_FF_3_net3512,
         cu0_RegisterBlock_FF_3_net3509, cu0_RegisterBlock_FF_3_net3500,
         cu0_RegisterBlock_1_FF_1_net3497, cu0_RegisterBlock_1_FF_1_net3494,
         cu1_counterChain_CounterRC_config__stride_0_,
         cu1_RegisterBlock_FF_1_net3506, cu1_RegisterBlock_FF_1_net3503,
         cu1_RegisterBlock_FF_1_net3500, cu1_RegisterBlock_FF_1_net3497,
         cu1_RegisterBlock_FF_1_net3494, cu1_RegisterBlock_FF_3_net3515,
         cu1_RegisterBlock_FF_3_net3512, cu1_RegisterBlock_FF_3_net3509,
         cu1_RegisterBlock_1_FF_1_net3518, cu1_RegisterBlock_1_FF_1_net3515,
         cu1_RegisterBlock_1_FF_1_net3497, cu1_RegisterBlock_1_FF_1_net3494,
         cu1_RegisterBlock_1_FF_1_net3491,
         cu1_controlBlock_UpDownCtr_1_reg__net3581,
         cu1_controlBlock_UpDownCtr_1_reg__net3578,
         cu1_controlBlock_UpDownCtr_1_reg__net3575,
         cu1_controlBlock_UpDownCtr_1_reg__net3572,
         cu0_controlBlock_UpDownCtr_reg__net3581,
         cu0_controlBlock_UpDownCtr_reg__net3578,
         cu0_controlBlock_UpDownCtr_reg__net3575,
         cu0_controlBlock_UpDownCtr_reg__net3572,
         cu0_controlBlock_UpDownCtr_1_reg__net3581,
         cu0_controlBlock_UpDownCtr_1_reg__net3578,
         cu0_controlBlock_UpDownCtr_1_reg__net3575,
         cu0_controlBlock_UpDownCtr_1_reg__net3572,
         cu1_controlBlock_UpDownCtr_reg__net3581,
         cu1_controlBlock_UpDownCtr_reg__net3578,
         cu1_controlBlock_UpDownCtr_reg__net3575,
         cu1_controlBlock_UpDownCtr_reg__net3572,
         cu0_counterChain_CounterRC_counter_reg__net3515,
         cu0_counterChain_CounterRC_counter_reg__net3512,
         cu0_counterChain_CounterRC_counter_reg__net3509,
         cu0_counterChain_CounterRC_1_counter_reg__net3515,
         cu0_counterChain_CounterRC_1_counter_reg__net3512,
         cu0_counterChain_CounterRC_1_counter_reg__net3509,
         cu1_counterChain_CounterRC_counter_reg__net3515,
         cu1_counterChain_CounterRC_counter_reg__net3512,
         cu1_counterChain_CounterRC_counter_reg__net3509,
         cu1_counterChain_CounterRC_1_counter_reg__net3518,
         cu1_counterChain_CounterRC_1_counter_reg__net3515,
         cu1_counterChain_CounterRC_1_counter_reg__net3512,
         cu1_counterChain_CounterRC_1_counter_reg__net3509, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416;
  wire   [2:0] cu1_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu1_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu1_RegisterBlock_io_passDataOut_2;
  wire   [2:0] cu0_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu0_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu0_RegisterBlock_io_passDataOut_2;
  wire   [6:5] cu0_RegisterBlock_io_passDataOut_3;
  wire   [5:3] cu1_IntFU_T7;
  wire   [2:0] cu0_mem0_mem;
  wire   [4:0] cu0_mem1_mem;
  wire   [4:3] cu0_IntFU_T7;
  wire   [7:0] cu1_mem0_mem;
  wire   [6:0] cu1_IntFU_1_m_T3;
  wire   [5:0] cu0_IntFU_1_m_T3;
  assign io_status = 1'b0;

  SNPS_CLOCK_GATE_HIGH_SRAM_0_33 cu0_mem1_clk_gate_mem_reg_0_ ( .CLK(clk), 
        .EN(cu0_mem0_N15), .ENCLK(cu0_mem1_net3732), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_32 cu0_mem1_clk_gate_mem_reg_1_ ( .CLK(clk), 
        .EN(cu0_mem0_N16), .ENCLK(cu0_mem1_net3727), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_31 cu0_mem1_clk_gate_mem_reg_2_ ( .CLK(clk), 
        .EN(cu0_mem0_N17), .ENCLK(cu0_mem1_net3722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_30 cu0_mem1_clk_gate_mem_reg_3_ ( .CLK(clk), 
        .EN(cu0_mem0_N18), .ENCLK(cu0_mem1_net3717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_29 cu0_mem1_clk_gate_mem_reg_4_ ( .CLK(clk), 
        .EN(cu0_mem0_N19), .ENCLK(cu0_mem1_net3712), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_28 cu0_mem1_clk_gate_mem_reg_5_ ( .CLK(clk), 
        .EN(cu0_mem0_N20), .ENCLK(cu0_mem1_net3707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_27 cu0_mem1_clk_gate_mem_reg_6_ ( .CLK(clk), 
        .EN(cu0_mem0_N21), .ENCLK(cu0_mem1_net3702), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_26 cu0_mem1_clk_gate_mem_reg_7_ ( .CLK(clk), 
        .EN(cu0_mem0_N22), .ENCLK(cu0_mem1_net3697), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_25 cu0_mem1_clk_gate_mem_reg_8_ ( .CLK(clk), 
        .EN(cu0_mem0_N23), .ENCLK(cu0_mem1_net3692), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_24 cu0_mem1_clk_gate_mem_reg_9_ ( .CLK(clk), 
        .EN(cu0_mem0_N24), .ENCLK(cu0_mem1_net3687), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_23 cu0_mem1_clk_gate_mem_reg_10_ ( .CLK(clk), 
        .EN(cu0_mem0_N25), .ENCLK(cu0_mem1_net3682), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_21 cu0_mem1_clk_gate_mem_reg_12_ ( .CLK(clk), 
        .EN(cu0_mem0_N27), .ENCLK(cu0_mem1_net3672), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_19 cu0_mem1_clk_gate_mem_reg_14_ ( .CLK(clk), 
        .EN(cu0_mem0_N29), .ENCLK(cu0_mem1_net3662), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_18 cu0_mem1_clk_gate_mem_reg_15_ ( .CLK(clk), 
        .EN(cu0_mem0_N30), .ENCLK(cu0_mem1_net3656), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_16 cu1_mem0_clk_gate_mem_reg_0_ ( .CLK(clk), 
        .EN(cu1_mem1_N15), .ENCLK(cu1_mem0_net3732), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_15 cu1_mem0_clk_gate_mem_reg_1_ ( .CLK(clk), 
        .EN(cu1_mem1_N16), .ENCLK(cu1_mem0_net3727), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_14 cu1_mem0_clk_gate_mem_reg_2_ ( .CLK(clk), 
        .EN(cu1_mem1_N17), .ENCLK(cu1_mem0_net3722), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_13 cu1_mem0_clk_gate_mem_reg_3_ ( .CLK(clk), 
        .EN(cu1_mem1_N18), .ENCLK(cu1_mem0_net3717), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_12 cu1_mem0_clk_gate_mem_reg_4_ ( .CLK(clk), 
        .EN(cu1_mem1_N19), .ENCLK(cu1_mem0_net3712), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_11 cu1_mem0_clk_gate_mem_reg_5_ ( .CLK(clk), 
        .EN(cu1_mem1_N20), .ENCLK(cu1_mem0_net3707), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_10 cu1_mem0_clk_gate_mem_reg_6_ ( .CLK(clk), 
        .EN(cu1_mem1_N21), .ENCLK(cu1_mem0_net3702), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_9 cu1_mem0_clk_gate_mem_reg_7_ ( .CLK(clk), .EN(
        cu1_mem1_N22), .ENCLK(cu1_mem0_net3697), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_8 cu1_mem0_clk_gate_mem_reg_8_ ( .CLK(clk), .EN(
        cu1_mem1_N23), .ENCLK(cu1_mem0_net3692), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_7 cu1_mem0_clk_gate_mem_reg_9_ ( .CLK(clk), .EN(
        cu1_mem1_N24), .ENCLK(cu1_mem0_net3687), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_6 cu1_mem0_clk_gate_mem_reg_10_ ( .CLK(clk), 
        .EN(cu1_mem1_N25), .ENCLK(cu1_mem0_net3682), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_4 cu1_mem0_clk_gate_mem_reg_12_ ( .CLK(clk), 
        .EN(cu1_mem1_N27), .ENCLK(cu1_mem0_net3672), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_2 cu1_mem0_clk_gate_mem_reg_14_ ( .CLK(clk), 
        .EN(cu1_mem1_N29), .ENCLK(cu1_mem0_net3662), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_SRAM_0_1 cu1_mem0_clk_gate_mem_reg_15_ ( .CLK(clk), 
        .EN(cu1_mem1_N30), .ENCLK(cu1_mem0_net3656), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 cu0_controlBlock_incXbar_clk_gate_config__outSelect_3_reg ( 
        .CLK(clk), .EN(cu0_controlBlock_incXbar_net3599), .ENCLK(
        cu0_controlBlock_incXbar_net3602), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_8 cu1_RegisterBlock_1_FF_1_clk_gate_ff_reg ( 
        .CLK(clk), .EN(cu1_RegisterBlock_1_FF_1_net3491), .ENCLK(
        cu1_RegisterBlock_1_FF_1_net3518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_1 cu1_counterChain_CounterRC_1_counter_reg__clk_gate_ff_reg ( 
        .CLK(clk), .EN(reset), .ENCLK(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .TE(1'b0) );
  DFQD4BWP cu1_mem1_mem_reg_1__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3727) );
  DFQD4BWP cu1_mem1_mem_reg_1__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3727) );
  DFQD4BWP cu1_mem1_mem_reg_1__7_ ( .D(n1416), .CP(cu1_mem0_net3727) );
  DFQD4BWP cu1_mem1_mem_reg_2__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3722) );
  DFQD4BWP cu1_mem1_mem_reg_2__6_ ( .D(n725), .CP(cu1_mem0_net3722) );
  DFQD4BWP cu1_mem1_mem_reg_2__7_ ( .D(n1416), .CP(cu1_mem0_net3722) );
  DFQD4BWP cu1_mem1_mem_reg_3__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3717) );
  DFQD4BWP cu1_mem1_mem_reg_3__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3717) );
  DFQD4BWP cu1_mem1_mem_reg_3__7_ ( .D(n1416), .CP(cu1_mem0_net3717) );
  DFQD4BWP cu1_mem1_mem_reg_4__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3712) );
  DFQD4BWP cu1_mem1_mem_reg_4__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3712) );
  DFQD4BWP cu1_mem1_mem_reg_4__7_ ( .D(n1416), .CP(cu1_mem0_net3712) );
  DFQD4BWP cu1_mem1_mem_reg_5__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3707) );
  DFQD4BWP cu1_mem1_mem_reg_5__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3707) );
  DFQD4BWP cu1_mem1_mem_reg_5__7_ ( .D(n1416), .CP(cu1_mem0_net3707) );
  DFQD4BWP cu1_mem1_mem_reg_6__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3702) );
  DFQD4BWP cu1_mem1_mem_reg_6__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3702) );
  DFQD4BWP cu1_mem1_mem_reg_6__7_ ( .D(n1416), .CP(cu1_mem0_net3702) );
  DFQD4BWP cu1_mem1_mem_reg_7__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3697) );
  DFQD4BWP cu1_mem1_mem_reg_7__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3697) );
  DFQD4BWP cu1_mem1_mem_reg_7__7_ ( .D(n1416), .CP(cu1_mem0_net3697) );
  DFQD4BWP cu1_mem1_mem_reg_8__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3692) );
  DFQD4BWP cu1_mem1_mem_reg_8__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3692) );
  DFQD4BWP cu1_mem1_mem_reg_8__7_ ( .D(n1416), .CP(cu1_mem0_net3692) );
  DFQD4BWP cu1_mem1_mem_reg_9__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3687) );
  DFQD4BWP cu1_mem1_mem_reg_9__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3687) );
  DFQD4BWP cu1_mem1_mem_reg_9__7_ ( .D(n1416), .CP(cu1_mem0_net3687) );
  DFQD4BWP cu1_mem1_mem_reg_10__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3682) );
  DFQD4BWP cu1_mem1_mem_reg_10__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3682) );
  DFQD4BWP cu1_mem1_mem_reg_10__7_ ( .D(n1416), .CP(cu1_mem0_net3682) );
  DFQD4BWP cu1_mem1_mem_reg_12__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3672) );
  DFQD4BWP cu1_mem1_mem_reg_12__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3672) );
  DFQD4BWP cu1_mem1_mem_reg_12__7_ ( .D(n1416), .CP(cu1_mem0_net3672) );
  DFQD4BWP cu1_mem1_mem_reg_14__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3662) );
  DFQD4BWP cu1_mem1_mem_reg_14__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3662) );
  DFQD4BWP cu1_mem1_mem_reg_14__7_ ( .D(n1416), .CP(cu1_mem0_net3662) );
  DFQD4BWP cu1_mem1_mem_reg_15__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3656) );
  DFQD4BWP cu1_mem1_mem_reg_15__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3656) );
  DFQD4BWP cu1_mem1_mem_reg_15__7_ ( .D(n1416), .CP(cu1_mem0_net3656) );
  DFQD4BWP cu1_controlBlock_config__udcInit_0_reg_1_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_mem0_mem_reg_1__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3727) );
  DFQD4BWP cu0_mem0_mem_reg_1__6_ ( .D(n1404), .CP(cu0_mem1_net3727) );
  DFQD4BWP cu0_mem0_mem_reg_1__7_ ( .D(n1405), .CP(cu0_mem1_net3727) );
  DFQD4BWP cu0_mem0_mem_reg_2__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3722) );
  DFQD4BWP cu0_mem0_mem_reg_2__6_ ( .D(n1404), .CP(cu0_mem1_net3722) );
  DFQD4BWP cu0_mem0_mem_reg_2__7_ ( .D(n1405), .CP(cu0_mem1_net3722) );
  DFQD4BWP cu0_mem0_mem_reg_3__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3717) );
  DFQD4BWP cu0_mem0_mem_reg_3__6_ ( .D(n1404), .CP(cu0_mem1_net3717) );
  DFQD4BWP cu0_mem0_mem_reg_3__7_ ( .D(n1405), .CP(cu0_mem1_net3717) );
  DFQD4BWP cu0_mem0_mem_reg_4__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3712) );
  DFQD4BWP cu0_mem0_mem_reg_4__6_ ( .D(n1404), .CP(cu0_mem1_net3712) );
  DFQD4BWP cu0_mem0_mem_reg_4__7_ ( .D(n1405), .CP(cu0_mem1_net3712) );
  DFQD4BWP cu0_mem0_mem_reg_5__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3707) );
  DFQD4BWP cu0_mem0_mem_reg_5__6_ ( .D(n1404), .CP(cu0_mem1_net3707) );
  DFQD4BWP cu0_mem0_mem_reg_5__7_ ( .D(n1405), .CP(cu0_mem1_net3707) );
  DFQD4BWP cu0_mem0_mem_reg_6__5_ ( .D(cu0_IntFU_1_m_T3[5]), .CP(
        cu0_mem1_net3702) );
  DFQD4BWP cu0_mem0_mem_reg_6__6_ ( .D(n1404), .CP(cu0_mem1_net3702) );
  DFQD4BWP cu0_mem0_mem_reg_6__7_ ( .D(n1405), .CP(cu0_mem1_net3702) );
  DFQD4BWP cu0_mem0_mem_reg_7__6_ ( .D(n1404), .CP(cu0_mem1_net3697) );
  DFQD4BWP cu0_mem0_mem_reg_7__7_ ( .D(n1405), .CP(cu0_mem1_net3697) );
  DFQD4BWP cu0_mem0_mem_reg_8__6_ ( .D(n1404), .CP(cu0_mem1_net3692) );
  DFQD4BWP cu0_mem0_mem_reg_8__7_ ( .D(n1405), .CP(cu0_mem1_net3692) );
  DFQD4BWP cu0_mem0_mem_reg_9__6_ ( .D(n1404), .CP(cu0_mem1_net3687) );
  DFQD4BWP cu0_mem0_mem_reg_9__7_ ( .D(n1405), .CP(cu0_mem1_net3687) );
  DFQD4BWP cu0_mem0_mem_reg_10__6_ ( .D(n1404), .CP(cu0_mem1_net3682) );
  DFQD4BWP cu0_mem0_mem_reg_10__7_ ( .D(n1405), .CP(cu0_mem1_net3682) );
  DFQD4BWP cu0_mem0_mem_reg_12__6_ ( .D(n1404), .CP(cu0_mem1_net3672) );
  DFQD4BWP cu0_mem0_mem_reg_12__7_ ( .D(n1405), .CP(cu0_mem1_net3672) );
  DFQD4BWP cu0_mem0_mem_reg_14__6_ ( .D(n1404), .CP(cu0_mem1_net3662) );
  DFQD4BWP cu0_mem0_mem_reg_14__7_ ( .D(n1405), .CP(cu0_mem1_net3662) );
  DFQD4BWP cu0_mem0_mem_reg_15__6_ ( .D(n1404), .CP(cu0_mem1_net3656) );
  DFQD4BWP cu0_mem0_mem_reg_15__7_ ( .D(n1405), .CP(cu0_mem1_net3656) );
  DFQD4BWP cu0_mem1_mem_reg_1__6_ ( .D(n1404), .CP(cu0_mem1_net3727) );
  DFQD4BWP cu0_mem1_mem_reg_1__7_ ( .D(n1405), .CP(cu0_mem1_net3727) );
  DFQD4BWP cu0_mem1_mem_reg_2__6_ ( .D(n1404), .CP(cu0_mem1_net3722) );
  DFQD4BWP cu0_mem1_mem_reg_2__7_ ( .D(n1405), .CP(cu0_mem1_net3722) );
  DFQD4BWP cu0_mem1_mem_reg_3__6_ ( .D(n1404), .CP(cu0_mem1_net3717) );
  DFQD4BWP cu0_mem1_mem_reg_3__7_ ( .D(n1405), .CP(cu0_mem1_net3717) );
  DFQD4BWP cu0_mem1_mem_reg_4__6_ ( .D(n1404), .CP(cu0_mem1_net3712) );
  DFQD4BWP cu0_mem1_mem_reg_4__7_ ( .D(n1405), .CP(cu0_mem1_net3712) );
  DFQD4BWP cu0_mem1_mem_reg_5__6_ ( .D(n1404), .CP(cu0_mem1_net3707) );
  DFQD4BWP cu0_mem1_mem_reg_5__7_ ( .D(n1405), .CP(cu0_mem1_net3707) );
  DFQD4BWP cu0_mem1_mem_reg_6__6_ ( .D(n1404), .CP(cu0_mem1_net3702) );
  DFQD4BWP cu0_mem1_mem_reg_6__7_ ( .D(n1405), .CP(cu0_mem1_net3702) );
  DFQD4BWP cu0_mem1_mem_reg_7__6_ ( .D(n1404), .CP(cu0_mem1_net3697) );
  DFQD4BWP cu0_mem1_mem_reg_7__7_ ( .D(n1405), .CP(cu0_mem1_net3697) );
  DFQD4BWP cu0_mem1_mem_reg_8__6_ ( .D(n1404), .CP(cu0_mem1_net3692) );
  DFQD4BWP cu0_mem1_mem_reg_8__7_ ( .D(n1405), .CP(cu0_mem1_net3692) );
  DFQD4BWP cu0_mem1_mem_reg_9__6_ ( .D(n1404), .CP(cu0_mem1_net3687) );
  DFQD4BWP cu0_mem1_mem_reg_9__7_ ( .D(n1405), .CP(cu0_mem1_net3687) );
  DFQD4BWP cu0_mem1_mem_reg_10__6_ ( .D(n1404), .CP(cu0_mem1_net3682) );
  DFQD4BWP cu0_mem1_mem_reg_10__7_ ( .D(n1405), .CP(cu0_mem1_net3682) );
  DFQD4BWP cu0_mem1_mem_reg_12__6_ ( .D(n1404), .CP(cu0_mem1_net3672) );
  DFQD4BWP cu0_mem1_mem_reg_12__7_ ( .D(n1405), .CP(cu0_mem1_net3672) );
  DFQD4BWP cu0_mem1_mem_reg_14__6_ ( .D(n1404), .CP(cu0_mem1_net3662) );
  DFQD4BWP cu0_mem1_mem_reg_14__7_ ( .D(n1405), .CP(cu0_mem1_net3662) );
  DFQD4BWP cu0_mem1_mem_reg_15__6_ ( .D(n1404), .CP(cu0_mem1_net3656) );
  DFQD4BWP cu0_mem1_mem_reg_15__7_ ( .D(n1405), .CP(cu0_mem1_net3656) );
  DFQD4BWP cu0_controlBlock_config__udcInit_0_reg_1_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu1_mem0_mem_reg_1__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3727) );
  DFQD4BWP cu1_mem0_mem_reg_1__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3727) );
  DFQD4BWP cu1_mem0_mem_reg_1__7_ ( .D(n1416), .CP(cu1_mem0_net3727) );
  DFQD4BWP cu1_mem0_mem_reg_2__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3722) );
  DFQD4BWP cu1_mem0_mem_reg_2__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3722) );
  DFQD4BWP cu1_mem0_mem_reg_2__7_ ( .D(n1416), .CP(cu1_mem0_net3722) );
  DFQD4BWP cu1_mem0_mem_reg_3__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3717) );
  DFQD4BWP cu1_mem0_mem_reg_3__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3717) );
  DFQD4BWP cu1_mem0_mem_reg_3__7_ ( .D(n1416), .CP(cu1_mem0_net3717) );
  DFQD4BWP cu1_mem0_mem_reg_4__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3712) );
  DFQD4BWP cu1_mem0_mem_reg_4__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3712) );
  DFQD4BWP cu1_mem0_mem_reg_4__7_ ( .D(n1416), .CP(cu1_mem0_net3712) );
  DFQD4BWP cu1_mem0_mem_reg_5__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3707) );
  DFQD4BWP cu1_mem0_mem_reg_5__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3707) );
  DFQD4BWP cu1_mem0_mem_reg_5__7_ ( .D(n1416), .CP(cu1_mem0_net3707) );
  DFQD4BWP cu1_mem0_mem_reg_6__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3702) );
  DFQD4BWP cu1_mem0_mem_reg_6__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3702) );
  DFQD4BWP cu1_mem0_mem_reg_6__7_ ( .D(n1416), .CP(cu1_mem0_net3702) );
  DFQD4BWP cu1_mem0_mem_reg_7__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3697) );
  DFQD4BWP cu1_mem0_mem_reg_7__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3697) );
  DFQD4BWP cu1_mem0_mem_reg_7__7_ ( .D(n1416), .CP(cu1_mem0_net3697) );
  DFQD4BWP cu1_mem0_mem_reg_8__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3692) );
  DFQD4BWP cu1_mem0_mem_reg_8__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3692) );
  DFQD4BWP cu1_mem0_mem_reg_8__7_ ( .D(n1416), .CP(cu1_mem0_net3692) );
  DFQD4BWP cu1_mem0_mem_reg_9__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3687) );
  DFQD4BWP cu1_mem0_mem_reg_9__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3687) );
  DFQD4BWP cu1_mem0_mem_reg_9__7_ ( .D(n1416), .CP(cu1_mem0_net3687) );
  DFQD4BWP cu1_mem0_mem_reg_10__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3682) );
  DFQD4BWP cu1_mem0_mem_reg_10__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3682) );
  DFQD4BWP cu1_mem0_mem_reg_10__7_ ( .D(n1416), .CP(cu1_mem0_net3682) );
  DFQD4BWP cu1_mem0_mem_reg_12__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3672) );
  DFQD4BWP cu1_mem0_mem_reg_12__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3672) );
  DFQD4BWP cu1_mem0_mem_reg_12__7_ ( .D(n1416), .CP(cu1_mem0_net3672) );
  DFQD4BWP cu1_mem0_mem_reg_14__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3662) );
  DFQD4BWP cu1_mem0_mem_reg_14__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3662) );
  DFQD4BWP cu1_mem0_mem_reg_14__7_ ( .D(n1416), .CP(cu1_mem0_net3662) );
  DFQD4BWP cu1_mem0_mem_reg_15__5_ ( .D(cu1_IntFU_1_m_T3[5]), .CP(
        cu1_mem0_net3656) );
  DFQD4BWP cu1_mem0_mem_reg_15__6_ ( .D(cu1_IntFU_1_m_T3[6]), .CP(
        cu1_mem0_net3656) );
  DFQD4BWP cu1_mem0_mem_reg_15__7_ ( .D(n1416), .CP(cu1_mem0_net3656) );
  DFQD4BWP cu1_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu1_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net3602) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_1_net3506), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_6_ ( .D(
        cu0_RegisterBlock_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_1_net3506), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_1_net3500), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_6_ ( .D(
        cu1_RegisterBlock_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_5_ ( .D(cu1_RegisterBlock_FF_1_net3500), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_6_ ( .D(cu0_RegisterBlock_FF_1_net3497), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_6_ ( .D(cu1_RegisterBlock_FF_1_net3497), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP controlBox_commandReg_reg ( .D(controlBox_N6), .CP(clk), .Q(
        controlBox_commandReg) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_7_ ( .D(cu1_RegisterBlock_FF_1_net3494), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD1BWP cu1_mem0_mem_reg_0__6_ ( .D(n725), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[6]) );
  DFQD1BWP cu1_mem0_mem_reg_0__7_ ( .D(n1416), .CP(cu1_mem0_net3732), .Q(
        cu1_mem0_mem[7]) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_5_ ( .D(cu0_RegisterBlock_FF_1_net3500), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_3_net3500), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[5]) );
  DFQD1BWP cu1_counterChain_CounterRC_config__stride_reg_0_ ( .D(reset), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_CounterRC_config__stride_0_) );
  DFQD2BWP cu1_RegisterBlock_1_FF_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3494), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD2BWP cu0_RegisterBlock_1_FF_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3494), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD2BWP cu0_RegisterBlock_FF_ff_reg_7_ ( .D(n731), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD2BWP cu0_RegisterBlock_FF_1_ff_reg_7_ ( .D(n731), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFQD1BWP cu1_RegisterBlock_FF_1_ff_reg_7_ ( .D(
        cu1_RegisterBlock_FF_1_net3494), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFD4BWP cu0_config__pipeStage_1_opB_value_reg_0_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net3602), .Q(n1403), .QN(n730) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_7_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_6_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_3_6_), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_5_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_4_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_3_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_2_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_1_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_0_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_7_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_6_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[6]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_5_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_4_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_3_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_2_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_1_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_4_ff_reg_0_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_2_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_0[2]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_1_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_0[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_2_ff_reg_0_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_0[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_7_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_6_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_3[6]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_5_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_3[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_4_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_3_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_2_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_1_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_5_ff_reg_0_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_7_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[7]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_6_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[6]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_5_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_4_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_3_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_2_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_1_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_4_ff_reg_0_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_2[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_2_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_0[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_1_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_0[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_2_ff_reg_0_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_0[0]), .CP(clk) );
  DFKCNQD1BWP controlBox_pulser_commandReg_reg ( .CN(n1415), .D(
        controlBox_commandReg), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_1_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[1]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_0_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[0]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_1_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[1]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_0_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[0]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_5_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[5]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_4_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[4]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_3_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[3]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_3_ff_reg_2_ ( .CN(n1415), .D(
        cu1_RegisterBlock_io_passDataOut_1[2]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_5_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[5]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_4_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[4]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_3_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[3]), .CP(clk) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_3_ff_reg_2_ ( .CN(n1415), .D(
        cu0_RegisterBlock_io_passDataOut_1[2]), .CP(clk) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_0_ ( .CN(n1411), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_0_ ( .CN(n1407), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_1_ ( .CN(n1412), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_1_ ( .CN(n1408), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem0_mem_reg_6__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem0_mem_reg_5__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem0_mem_reg_4__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem0_mem_reg_3__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem0_mem_reg_2__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem0_mem_reg_1__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu1_mem1_mem_reg_15__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem1_mem_reg_14__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem1_mem_reg_12__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem1_mem_reg_10__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem1_mem_reg_9__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem1_mem_reg_8__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem1_mem_reg_7__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem1_mem_reg_6__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem1_mem_reg_5__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem1_mem_reg_4__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem1_mem_reg_3__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem1_mem_reg_2__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem1_mem_reg_1__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu1_mem0_mem_reg_15__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3656) );
  DFKCNQD1BWP cu1_mem0_mem_reg_14__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3662) );
  DFKCNQD1BWP cu1_mem0_mem_reg_12__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3672) );
  DFKCNQD1BWP cu1_mem0_mem_reg_10__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3682) );
  DFKCNQD1BWP cu1_mem0_mem_reg_9__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3687) );
  DFKCNQD1BWP cu1_mem0_mem_reg_8__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3692) );
  DFKCNQD1BWP cu1_mem0_mem_reg_7__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3697) );
  DFKCNQD1BWP cu1_mem0_mem_reg_6__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3702) );
  DFKCNQD1BWP cu1_mem0_mem_reg_5__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3707) );
  DFKCNQD1BWP cu1_mem0_mem_reg_4__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3712) );
  DFKCNQD1BWP cu1_mem0_mem_reg_3__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3717) );
  DFKCNQD1BWP cu1_mem0_mem_reg_2__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3722) );
  DFKCNQD1BWP cu1_mem0_mem_reg_1__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3727) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_1_ff_reg_2_ ( .CN(n1413), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_1_ff_reg_2_ ( .CN(n1409), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518) );
  DFKCNQD1BWP cu0_mem1_mem_reg_15__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem1_mem_reg_14__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem1_mem_reg_12__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem1_mem_reg_10__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem1_mem_reg_9__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem1_mem_reg_8__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem1_mem_reg_7__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu0_mem1_mem_reg_6__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3702) );
  DFKCNQD1BWP cu0_mem1_mem_reg_5__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3707) );
  DFKCNQD1BWP cu0_mem1_mem_reg_4__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3712) );
  DFKCNQD1BWP cu0_mem1_mem_reg_3__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3717) );
  DFKCNQD1BWP cu0_mem1_mem_reg_2__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3722) );
  DFKCNQD1BWP cu0_mem1_mem_reg_1__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3727) );
  DFKCNQD1BWP cu0_mem0_mem_reg_15__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3656) );
  DFKCNQD1BWP cu0_mem0_mem_reg_14__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3662) );
  DFKCNQD1BWP cu0_mem0_mem_reg_12__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3672) );
  DFKCNQD1BWP cu0_mem0_mem_reg_10__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3682) );
  DFKCNQD1BWP cu0_mem0_mem_reg_9__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3687) );
  DFKCNQD1BWP cu0_mem0_mem_reg_8__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3692) );
  DFKCNQD1BWP cu0_mem0_mem_reg_7__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3697) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_5_ff_reg_6_ ( .CN(n1415), .D(
        cu1_mem1_mem_0__6_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3_6_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_6_ ( .CN(n1415), .D(
        cu1_mem0_mem[6]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[6])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_5_ff_reg_6_ ( .CN(n1415), .D(
        cu0_mem0_mem[1]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_3[6])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_5_ff_reg_5_ ( .CN(n1415), .D(
        cu0_mem0_mem[0]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_3[5])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_6_ ( .CN(n1415), .D(
        cu0_mem0_mem[1]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[6])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_5_ ( .CN(n1415), .D(
        cu0_mem0_mem[0]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[5])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_7_ ( .CN(n1415), .D(
        cu0_mem0_mem[2]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[7])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_7_ ( .CN(n1415), .D(
        cu1_mem0_mem[7]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[7])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_5_ ( .CN(n1415), .D(
        cu1_mem0_mem[5]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[5])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_4_ ( .CN(n1415), .D(
        cu1_mem0_mem[4]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[4])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_3_ ( .CN(n1415), .D(
        cu1_mem0_mem[3]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[3])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_2_ ( .CN(n1415), .D(
        cu1_mem0_mem[2]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[2])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_1_ ( .CN(n1415), .D(
        cu1_mem0_mem[1]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[1])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_4_ff_reg_0_ ( .CN(n1415), .D(
        cu1_mem0_mem[0]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_2[0])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_4_ ( .CN(n1415), .D(
        cu0_mem1_mem[4]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[4])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_3_ ( .CN(n1415), .D(
        cu0_mem1_mem[3]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[3])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_2_ ( .CN(n1415), .D(
        cu0_mem1_mem[2]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[2])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_1_ ( .CN(n1415), .D(
        cu0_mem1_mem[1]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[1])
         );
  DFKCNQD1BWP cu0_RegisterBlock_FF_4_ff_reg_0_ ( .CN(n1415), .D(
        cu0_mem1_mem[0]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_2[0])
         );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_2_ ( .CN(n1415), .D(
        cu1_counterChain_io_data_0_out_2_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[2]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_2_ ( .CN(n1415), .D(
        cu0_counterChain_io_data_0_out_2_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[2]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_1_ ( .CN(n1415), .D(
        cu0_counterChain_io_data_0_out_1_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[1]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_1_ ( .CN(n1415), .D(
        cu1_counterChain_io_data_0_out_1_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[1]) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3581), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_2_ff_reg_0_ ( .CN(n1415), .D(
        cu0_counterChain_io_data_0_out_0_), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[0]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_0_ ( .CN(n1415), .D(
        cu1_counterChain_io_data_0_out_0_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[0]) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_0_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_0_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_2_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_0_out_1_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_2_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_0_out_1_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_1_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_0_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3515), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_0_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_1_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_2_) );
  DFKCNQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu0_counterChain_CounterRC_1_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_counterChain_io_data_1_out_1_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3509), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_2_) );
  DFKCNQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .CN(1'b1), 
        .D(cu1_counterChain_CounterRC_1_counter_reg__net3512), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_counterChain_io_data_1_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3578), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3575), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_1_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFKCNQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu1_controlBlock_UpDownCtr_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_1_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFKCNQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .CN(1'b1), .D(
        cu0_controlBlock_UpDownCtr_reg__net3572), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_0_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_3_net3515), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[0]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_3_ff_reg_0_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_3_net3515), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[0]) );
  DFKCNQD1BWP cu0_mem1_mem_reg_0__0_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[0]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem1_mem[0]) );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__0_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[0]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[0]) );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__1_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[1]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[1]) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_0_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[0]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_0_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[0]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_0_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_3_ff_reg_1_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_3_net3512), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[1]) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_0_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_1_FF_1_net3515), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_0_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[0]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_0_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_0_ ( .CN(n1411), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_0_) );
  DFKCNQD1BWP cu0_mem1_mem_reg_0__1_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[1]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem1_mem[1]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_1_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_3_net3512), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[1]) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_1_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[1]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_1_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[1]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_1_) );
  DFKCNQD1BWP cu0_mem1_mem_reg_0__2_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[2]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem1_mem[2]) );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__2_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[2]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[2]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_0_ ( .CN(n1407), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_0_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_1_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[1]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_1_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[1]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_1_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_1_ ( .CN(n1412), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_1_) );
  DFKCNQD1BWP cu0_mem1_mem_reg_0__3_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[3]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem1_mem[3]) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_2_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[2]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_2_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[2]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_2_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_1_ ( .CN(n1408), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_1_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_2_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[2]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_2_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[2]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_2_) );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__3_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[3]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[3]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_3_ff_reg_2_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_3_net3509), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[2]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_2_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_3_net3509), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[2]) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_3_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[3]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_3_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[3]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_3_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_3_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[3]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_3_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[3]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_3_) );
  DFKCNQD1BWP cu0_mem1_mem_reg_0__4_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[4]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem1_mem[4]) );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__4_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[4]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[4]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_3_ff_reg_3_ ( .CN(cu0_IntFU_T7[3]), .D(
        n1406), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_1[3]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_3_ ( .CN(cu1_IntFU_T7[3]), .D(
        n1406), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_1[3]) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_2_ ( .CN(n1413), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_2_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_2_ ( .CN(n1409), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_2_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_4_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[4]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_4_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[4]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_4_) );
  DFKCNQD1BWP cu0_mem0_mem_reg_0__5_ ( .CN(1'b1), .D(cu0_IntFU_1_m_T3[5]), 
        .CP(cu0_mem1_net3732), .Q(cu0_mem0_mem[0]) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_4_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[4]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_4_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[4]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_4_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_4_ ( .CN(n1406), .D(
        cu1_IntFU_T7[4]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_1[4])
         );
  DFKCNQD1BWP cu1_mem0_mem_reg_0__5_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[5]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem0_mem[5]) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_4_ ( .CN(1'b1), .D(
        cu1_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_4_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_3_ ( .CN(n1414), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_3_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_3_ff_reg_4_ ( .CN(n1406), .D(
        cu0_IntFU_T7[4]), .CP(clk), .Q(cu0_RegisterBlock_io_passDataOut_1[4])
         );
  DFKCNQD1BWP cu1_mem1_mem_reg_0__6_ ( .CN(1'b1), .D(cu1_IntFU_1_m_T3[6]), 
        .CP(cu1_mem0_net3732), .Q(cu1_mem1_mem_0__6_) );
  DFKCNQD1BWP cu0_RegisterBlock_FF_ff_reg_4_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_FF_1_net3503), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_FF_io_data_out_4_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_ff_reg_3_ ( .CN(n728), .D(n1415), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_FF_io_data_out_3_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_5_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[5]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_5_ ( .CN(n1415), .D(
        cu0_IntFU_1_m_T3[5]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_5_) );
  DFKCNQD1BWP cu0_mem0_mem_reg_0__6_ ( .CN(1'b1), .D(n1404), .CP(
        cu0_mem1_net3732), .Q(cu0_mem0_mem[1]) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_6_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFKCNQD1BWP cu0_RegisterBlock_1_FF_ff_reg_6_ ( .CN(1'b1), .D(
        cu0_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_6_) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_3_ff_reg_5_ ( .CN(n1406), .D(
        cu1_IntFU_T7[5]), .CP(clk), .Q(cu1_RegisterBlock_io_passDataOut_1[5])
         );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_5_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[5]), .CP(cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_ff_reg_5_ ( .CN(n1415), .D(
        cu1_IntFU_1_m_T3[5]), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3494), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_7_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_1_net3494), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_7_) );
  DFQD1BWP cu0_mem0_mem_reg_0__7_ ( .D(n1405), .CP(cu0_mem1_net3732), .Q(
        cu0_mem0_mem[2]) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net3518), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net3497), .CP(
        cu1_RegisterBlock_1_FF_1_net3518), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFQD4BWP cu1_mem0_mem_reg_13__6_ ( .D(n712), .CP(clk), .Q(n712) );
  DFQD4BWP cu1_mem0_mem_reg_13__7_ ( .D(n711), .CP(clk), .Q(n711) );
  DFQD4BWP cu1_mem1_mem_reg_13__7_ ( .D(n710), .CP(clk), .Q(n710) );
  DFQD4BWP cu1_mem1_mem_reg_13__6_ ( .D(n709), .CP(clk), .Q(n709) );
  DFQD4BWP cu1_mem1_mem_reg_13__0_ ( .D(n708), .CP(clk), .Q(n708) );
  DFQD4BWP cu1_mem0_mem_reg_13__0_ ( .D(n707), .CP(clk), .Q(n707) );
  DFQD4BWP cu1_mem1_mem_reg_13__1_ ( .D(n706), .CP(clk), .Q(n706) );
  DFQD4BWP cu1_mem0_mem_reg_13__1_ ( .D(n705), .CP(clk), .Q(n705) );
  DFQD4BWP cu1_mem1_mem_reg_13__2_ ( .D(n704), .CP(clk), .Q(n704) );
  DFQD4BWP cu1_mem0_mem_reg_13__2_ ( .D(n703), .CP(clk), .Q(n703) );
  DFQD4BWP cu1_mem1_mem_reg_13__3_ ( .D(n702), .CP(clk), .Q(n702) );
  DFQD4BWP cu1_mem0_mem_reg_13__3_ ( .D(n701), .CP(clk), .Q(n701) );
  DFQD4BWP cu1_mem1_mem_reg_13__4_ ( .D(n700), .CP(clk), .Q(n700) );
  DFQD4BWP cu1_mem0_mem_reg_13__4_ ( .D(n699), .CP(clk), .Q(n699) );
  DFQD4BWP cu1_mem0_mem_reg_13__5_ ( .D(n698), .CP(clk), .Q(n698) );
  DFQD4BWP cu1_mem1_mem_reg_13__5_ ( .D(n697), .CP(clk), .Q(n697) );
  DFQD4BWP cu0_mem1_mem_reg_11__6_ ( .D(n696), .CP(clk), .Q(n696) );
  DFQD4BWP cu0_mem0_mem_reg_11__5_ ( .D(n695), .CP(clk), .Q(n695) );
  DFQD4BWP cu0_mem1_mem_reg_11__5_ ( .D(n694), .CP(clk), .Q(n694) );
  DFQD4BWP cu0_mem0_mem_reg_11__4_ ( .D(n693), .CP(clk), .Q(n693) );
  DFQD4BWP cu0_mem1_mem_reg_11__4_ ( .D(n692), .CP(clk), .Q(n692) );
  DFQD4BWP cu0_mem0_mem_reg_11__3_ ( .D(n691), .CP(clk), .Q(n691) );
  DFQD4BWP cu0_mem1_mem_reg_11__3_ ( .D(n690), .CP(clk), .Q(n690) );
  DFQD4BWP cu0_mem0_mem_reg_11__2_ ( .D(n689), .CP(clk), .Q(n689) );
  DFQD4BWP cu0_mem1_mem_reg_11__2_ ( .D(n688), .CP(clk), .Q(n688) );
  DFQD4BWP cu0_mem0_mem_reg_11__1_ ( .D(n687), .CP(clk), .Q(n687) );
  DFQD4BWP cu0_mem1_mem_reg_11__1_ ( .D(n686), .CP(clk), .Q(n686) );
  DFQD4BWP cu0_mem0_mem_reg_11__0_ ( .D(n685), .CP(clk), .Q(n685) );
  DFQD4BWP cu0_mem1_mem_reg_11__0_ ( .D(n684), .CP(clk), .Q(n684) );
  DFQD4BWP cu0_mem0_mem_reg_11__6_ ( .D(n683), .CP(clk), .Q(n683) );
  DFQD4BWP cu0_mem0_mem_reg_11__7_ ( .D(n682), .CP(clk), .Q(n682) );
  DFQD4BWP cu0_mem1_mem_reg_11__7_ ( .D(n681), .CP(clk), .Q(n681) );
  DFQD4BWP cu0_mem1_mem_reg_13__6_ ( .D(n680), .CP(clk), .Q(n680) );
  DFQD4BWP cu0_mem0_mem_reg_13__5_ ( .D(n679), .CP(clk), .Q(n679) );
  DFQD4BWP cu0_mem1_mem_reg_13__5_ ( .D(n678), .CP(clk), .Q(n678) );
  DFQD4BWP cu0_mem0_mem_reg_13__4_ ( .D(n677), .CP(clk), .Q(n677) );
  DFQD4BWP cu0_mem1_mem_reg_13__4_ ( .D(n676), .CP(clk), .Q(n676) );
  DFQD4BWP cu0_mem0_mem_reg_13__3_ ( .D(n675), .CP(clk), .Q(n675) );
  DFQD4BWP cu0_mem1_mem_reg_13__3_ ( .D(n674), .CP(clk), .Q(n674) );
  DFQD4BWP cu0_mem0_mem_reg_13__2_ ( .D(n673), .CP(clk), .Q(n673) );
  DFQD4BWP cu0_mem1_mem_reg_13__2_ ( .D(n672), .CP(clk), .Q(n672) );
  DFQD4BWP cu0_mem0_mem_reg_13__1_ ( .D(n671), .CP(clk), .Q(n671) );
  DFQD4BWP cu0_mem1_mem_reg_13__1_ ( .D(n670), .CP(clk), .Q(n670) );
  DFQD4BWP cu0_mem0_mem_reg_13__0_ ( .D(n669), .CP(clk), .Q(n669) );
  DFQD4BWP cu0_mem1_mem_reg_13__0_ ( .D(n668), .CP(clk), .Q(n668) );
  DFQD4BWP cu0_mem0_mem_reg_13__6_ ( .D(n667), .CP(clk), .Q(n667) );
  DFQD4BWP cu0_mem0_mem_reg_13__7_ ( .D(n666), .CP(clk), .Q(n666) );
  DFQD4BWP cu0_mem1_mem_reg_13__7_ ( .D(n665), .CP(clk), .Q(n665) );
  DFQD4BWP cu1_mem1_mem_reg_11__5_ ( .D(n664), .CP(clk), .Q(n664) );
  DFQD4BWP cu1_mem0_mem_reg_11__5_ ( .D(n663), .CP(clk), .Q(n663) );
  DFQD4BWP cu1_mem0_mem_reg_11__4_ ( .D(n662), .CP(clk), .Q(n662) );
  DFQD4BWP cu1_mem1_mem_reg_11__4_ ( .D(n661), .CP(clk), .Q(n661) );
  DFQD4BWP cu1_mem0_mem_reg_11__3_ ( .D(n660), .CP(clk), .Q(n660) );
  DFQD4BWP cu1_mem1_mem_reg_11__3_ ( .D(n659), .CP(clk), .Q(n659) );
  DFQD4BWP cu1_mem0_mem_reg_11__2_ ( .D(n658), .CP(clk), .Q(n658) );
  DFQD4BWP cu1_mem1_mem_reg_11__2_ ( .D(n657), .CP(clk), .Q(n657) );
  DFQD4BWP cu1_mem0_mem_reg_11__1_ ( .D(n656), .CP(clk), .Q(n656) );
  DFQD4BWP cu1_mem1_mem_reg_11__1_ ( .D(n655), .CP(clk), .Q(n655) );
  DFQD4BWP cu1_mem0_mem_reg_11__0_ ( .D(n654), .CP(clk), .Q(n654) );
  DFQD4BWP cu1_mem1_mem_reg_11__0_ ( .D(n653), .CP(clk), .Q(n653) );
  DFQD4BWP cu1_mem1_mem_reg_11__6_ ( .D(n652), .CP(clk), .Q(n652) );
  DFQD4BWP cu1_mem1_mem_reg_11__7_ ( .D(n651), .CP(clk), .Q(n651) );
  DFQD4BWP cu1_mem0_mem_reg_11__7_ ( .D(n650), .CP(clk), .Q(n650) );
  DFQD4BWP cu1_mem0_mem_reg_11__6_ ( .D(n649), .CP(clk), .Q(n649) );
  FICIND2BWP U972 ( .CIN(n761), .B(1'b0), .A(n763), .S(n764) );
  INVD1BWP U973 ( .I(n833), .ZN(n864) );
  INVD1BWP U974 ( .I(n995), .ZN(n942) );
  INVD1BWP U975 ( .I(n840), .ZN(n930) );
  INVD1BWP U976 ( .I(n816), .ZN(n932) );
  INVD1BWP U977 ( .I(n730), .ZN(n726) );
  INVD1BWP U978 ( .I(n883), .ZN(n863) );
  INVD1BWP U979 ( .I(n826), .ZN(n862) );
  ND2D1BWP U980 ( .A1(n730), .A2(cu0_RegisterBlock_FF_io_data_out_2_), .ZN(
        n736) );
  INVD1BWP U981 ( .I(n834), .ZN(n860) );
  INVD1BWP U982 ( .I(n929), .ZN(n938) );
  INVD1BWP U983 ( .I(n817), .ZN(n941) );
  FA1D1BWP U984 ( .A(n919), .B(n918), .CI(n917), .CO(n920), .S(n786) );
  IOA21D1BWP U985 ( .A1(cu1_counterChain_io_data_1_out_2_), .A2(n1403), .B(
        n778), .ZN(n817) );
  ND2D1BWP U986 ( .A1(n778), .A2(n772), .ZN(n816) );
  IOA21D1BWP U987 ( .A1(n1403), .A2(cu0_counterChain_io_data_1_out_2_), .B(
        n736), .ZN(n825) );
  IOA21D1BWP U988 ( .A1(n1403), .A2(cu0_counterChain_io_data_0_out_2_), .B(
        n736), .ZN(n826) );
  IND2D1BWP U989 ( .A1(n781), .B1(n780), .ZN(n839) );
  INR2D1BWP U990 ( .A1(n1403), .B1(n779), .ZN(n781) );
  ND2D1BWP U991 ( .A1(n780), .A2(n774), .ZN(n840) );
  IND2D1BWP U992 ( .A1(n740), .B1(n739), .ZN(n833) );
  IND2D1BWP U993 ( .A1(n740), .B1(n737), .ZN(n834) );
  ND2D1BWP U994 ( .A1(n1403), .A2(cu0_counterChain_io_data_1_out_1_), .ZN(n737) );
  ND2D1BWP U995 ( .A1(n729), .A2(n742), .ZN(n824) );
  NR2D1BWP U996 ( .A1(n776), .A2(n784), .ZN(n937) );
  NR2D1BWP U997 ( .A1(n730), .A2(n783), .ZN(n784) );
  INVD1BWP U998 ( .I(n824), .ZN(n846) );
  INVD1BWP U999 ( .I(n827), .ZN(n845) );
  AN2XD1BWP U1000 ( .A1(n730), .A2(cu0_RegisterBlock_FF_io_data_out_3_), .Z(
        n883) );
  OAI22D1BWP U1001 ( .A1(n727), .A2(n760), .B1(n766), .B2(n765), .ZN(n761) );
  IOA21D1BWP U1002 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_6_), 
        .B(n759), .ZN(n765) );
  INVD1BWP U1003 ( .I(n759), .ZN(n766) );
  OR2XD1BWP U1004 ( .A1(n1414), .A2(n1413), .Z(n978) );
  INR2D1BWP U1005 ( .A1(n1413), .B1(n1414), .ZN(n975) );
  INVD1BWP U1006 ( .I(n948), .ZN(n734) );
  INVD1BWP U1007 ( .I(n949), .ZN(n735) );
  NR2D1BWP U1008 ( .A1(n786), .A2(n785), .ZN(n924) );
  ND2D1BWP U1009 ( .A1(n730), .A2(cu1_RegisterBlock_1_FF_io_data_out_4_), .ZN(
        n748) );
  OAI22D1BWP U1010 ( .A1(n810), .A2(n809), .B1(n808), .B2(n807), .ZN(n894) );
  NR2D1BWP U1011 ( .A1(n879), .A2(n878), .ZN(n880) );
  INVD1BWP U1012 ( .I(n955), .ZN(n879) );
  INR2D1BWP U1013 ( .A1(n1415), .B1(n726), .ZN(n996) );
  INR2D1BWP U1014 ( .A1(n726), .B1(reset), .ZN(n1406) );
  HICOND1BWP U1015 ( .A(n889), .CI(n888), .CON(n906), .S(cu1_IntFU_1_m_T3[0])
         );
  IOA21D1BWP U1016 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_0_), 
        .B(n758), .ZN(n889) );
  INR2D1BWP U1017 ( .A1(n1415), .B1(n887), .ZN(
        cu1_RegisterBlock_1_FF_1_net3494) );
  IOA21D1BWP U1018 ( .A1(n1403), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_5_), 
        .B(n797), .ZN(n892) );
  IOA21D1BWP U1019 ( .A1(n1403), .A2(cu0_counterChain_io_data_1_out_0_), .B(
        n729), .ZN(n827) );
  IND2D1BWP U1020 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_1_), 
        .ZN(n769) );
  IND2D1BWP U1021 ( .A1(n1413), .B1(n1414), .ZN(n974) );
  AN2XD1BWP U1022 ( .A1(n940), .A2(n939), .Z(n944) );
  XOR3D1BWP U1023 ( .A1(n935), .A2(n934), .A3(n933), .Z(n946) );
  XOR3D1BWP U1024 ( .A1(n947), .A2(n946), .A3(n945), .Z(n950) );
  CKND1BWP U1025 ( .I(n726), .ZN(n713) );
  AN3D1BWP U1026 ( .A1(n713), .A2(n996), .A3(
        cu1_RegisterBlock_FF_io_data_out_6_), .Z(
        cu1_RegisterBlock_FF_1_net3494) );
  NR2D1BWP U1027 ( .A1(n861), .A2(n864), .ZN(n714) );
  NR2D1BWP U1028 ( .A1(n863), .A2(n845), .ZN(n715) );
  CKXOR2D1BWP U1029 ( .A1(n714), .A2(n715), .Z(n849) );
  AN2D1BWP U1030 ( .A1(n714), .A2(n715), .Z(n869) );
  IND2D1BWP U1031 ( .A1(n1412), .B1(n973), .ZN(n979) );
  IND2D1BWP U1032 ( .A1(n1408), .B1(n1407), .ZN(n990) );
  OR2D1BWP U1033 ( .A1(n921), .A2(n920), .Z(n952) );
  IND3D1BWP U1034 ( .A1(cu1_counterChain_io_data_1_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n1415), .ZN(n1024)
         );
  IOA21D1BWP U1035 ( .A1(n1403), .A2(cu0_RegisterBlock_io_passDataOut_1[1]), 
        .B(n769), .ZN(n805) );
  AN3D1BWP U1036 ( .A1(n716), .A2(n996), .A3(
        cu1_RegisterBlock_FF_io_data_out_5_), .Z(
        cu1_RegisterBlock_FF_1_net3497) );
  CKND1BWP U1037 ( .I(n726), .ZN(n716) );
  IND2D1BWP U1038 ( .A1(n1408), .B1(n984), .ZN(n993) );
  IND3D1BWP U1039 ( .A1(cu0_counterChain_io_data_1_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n1415), .ZN(n1020)
         );
  ND2D1BWP U1040 ( .A1(n827), .A2(n824), .ZN(n832) );
  IND2D1BWP U1041 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_2_), 
        .ZN(n803) );
  IOA21D1BWP U1042 ( .A1(n1403), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_1_), 
        .B(n769), .ZN(n806) );
  AO22D1BWP U1043 ( .A1(n996), .A2(n929), .B1(n1406), .B2(cu1_IntFU_T7[5]), 
        .Z(cu1_RegisterBlock_FF_1_net3500) );
  NR2D1BWP U1044 ( .A1(n849), .A2(n850), .ZN(n876) );
  IND3D1BWP U1045 ( .A1(cu0_counterChain_io_data_0_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n1415), .ZN(n1018)
         );
  OA21D1BWP U1046 ( .A1(n843), .A2(n842), .B(n844), .Z(n965) );
  OA21D1BWP U1047 ( .A1(n837), .A2(n836), .B(n838), .Z(n964) );
  INR2D1BWP U1048 ( .A1(cu0_RegisterBlock_FF_io_data_out_4_), .B1(n1403), .ZN(
        n970) );
  AN2D1BWP U1049 ( .A1(n730), .A2(cu0_RegisterBlock_FF_io_data_out_5_), .Z(
        n743) );
  AO21D1BWP U1050 ( .A1(n730), .A2(n822), .B(n966), .Z(n1409) );
  AO21D1BWP U1051 ( .A1(n730), .A2(n831), .B(n967), .Z(n1413) );
  AOI21D1BWP U1052 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_3_), .A2(n1403), 
        .B(n717), .ZN(n718) );
  IAO21D1BWP U1053 ( .A1(n730), .A2(n802), .B(n717), .ZN(n719) );
  XNR3D1BWP U1054 ( .A1(n893), .A2(n718), .A3(n719), .ZN(cu0_IntFU_1_m_T3[3])
         );
  MAOI222D1BWP U1055 ( .A(n893), .B(n718), .C(n719), .ZN(n897) );
  CKND1BWP U1056 ( .I(n801), .ZN(n717) );
  XNR3D1BWP U1057 ( .A1(n805), .A2(n810), .A3(n806), .ZN(cu0_IntFU_1_m_T3[1])
         );
  AO22D1BWP U1058 ( .A1(n996), .A2(n995), .B1(n1406), .B2(cu1_IntFU_T7[4]), 
        .Z(cu1_RegisterBlock_FF_1_net3503) );
  IND2D1BWP U1059 ( .A1(n1403), .B1(cu1_RegisterBlock_FF_io_data_out_2_), .ZN(
        n778) );
  AO21D1BWP U1060 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_6_), .A2(n1403), 
        .B(n811), .Z(n857) );
  IND3D1BWP U1061 ( .A1(cu1_counterChain_io_data_0_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n1415), .ZN(n1022)
         );
  IND2D1BWP U1062 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_4_), 
        .ZN(n799) );
  IND2D1BWP U1063 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_3_), 
        .ZN(n801) );
  IND2D1BWP U1064 ( .A1(n1403), .B1(cu1_RegisterBlock_1_FF_io_data_out_2_), 
        .ZN(n752) );
  IND2D1BWP U1065 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_5_), 
        .ZN(n797) );
  INR2D1BWP U1066 ( .A1(n725), .B1(reset), .ZN(
        cu1_RegisterBlock_1_FF_1_net3497) );
  NR2D1BWP U1067 ( .A1(n734), .A2(n735), .ZN(n720) );
  IOA21D1BWP U1068 ( .A1(n953), .A2(n952), .B(n951), .ZN(n721) );
  XOR3D1BWP U1069 ( .A1(n720), .A2(n950), .A3(n721), .Z(cu1_IntFU_T7[5]) );
  INR2D1BWP U1070 ( .A1(cu1_IntFU_1_m_T3[0]), .B1(reset), .ZN(
        cu1_RegisterBlock_1_FF_1_net3515) );
  AO21D1BWP U1071 ( .A1(n841), .A2(n730), .B(n965), .Z(n1408) );
  AO21D1BWP U1072 ( .A1(n835), .A2(n730), .B(n964), .Z(n1412) );
  IOA21D1BWP U1073 ( .A1(n1403), .A2(cu0_RegisterBlock_io_passDataOut_1[0]), 
        .B(n771), .ZN(n722) );
  CKND2D1BWP U1074 ( .A1(n771), .A2(n770), .ZN(n723) );
  CKND2D1BWP U1075 ( .A1(n722), .A2(n723), .ZN(n810) );
  CKXOR2D1BWP U1076 ( .A1(n722), .A2(n723), .Z(cu0_IntFU_1_m_T3[0]) );
  AO22D1BWP U1077 ( .A1(n996), .A2(n997), .B1(n1406), .B2(cu0_IntFU_T7[4]), 
        .Z(cu0_RegisterBlock_FF_1_net3503) );
  INR2D1BWP U1078 ( .A1(n1414), .B1(reset), .ZN(cu0_RegisterBlock_FF_1_net3506) );
  CKND2D2BWP U1079 ( .A1(cu1_RegisterBlock_1_FF_io_data_out_1_), .A2(n730), 
        .ZN(n724) );
  XOR2D1BWP U1080 ( .A1(n768), .A2(n767), .Z(n725) );
  XOR2D2BWP U1081 ( .A1(n768), .A2(n767), .Z(cu1_IntFU_1_m_T3[6]) );
  FICIND2BWP U1082 ( .CIN(n900), .B(n901), .A(n902), .CO(n727) );
  CKAN2D1BWP U1083 ( .A1(n1403), .A2(cu1_counterChain_io_data_0_out_0_), .Z(
        n777) );
  CKND2D3BWP U1084 ( .A1(n886), .A2(n885), .ZN(n1414) );
  CKND2BWP U1085 ( .I(n983), .ZN(n985) );
  XOR2D2BWP U1086 ( .A1(n814), .A2(n813), .Z(n732) );
  CKND2BWP U1087 ( .I(n986), .ZN(n987) );
  INR2D2BWP U1088 ( .A1(n989), .B1(n1410), .ZN(n986) );
  INVD1BWP U1089 ( .I(n971), .ZN(n728) );
  CKND2D3BWP U1090 ( .A1(n796), .A2(n795), .ZN(n1410) );
  OR2XD1BWP U1091 ( .A1(n1403), .A2(n741), .Z(n729) );
  AN2XD1BWP U1092 ( .A1(n745), .A2(n996), .Z(n731) );
  INR2D1BWP U1093 ( .A1(cu0_RegisterBlock_1_FF_io_data_out_6_), .B1(n1403), 
        .ZN(n811) );
  INVD1BWP U1094 ( .I(n776), .ZN(n782) );
  NR2D1BWP U1095 ( .A1(n1403), .A2(n775), .ZN(n776) );
  INR2D1BWP U1096 ( .A1(cu1_RegisterBlock_FF_io_data_out_4_), .B1(n1403), .ZN(
        n929) );
  INR2D1BWP U1097 ( .A1(n782), .B1(n777), .ZN(n936) );
  OR2XD1BWP U1098 ( .A1(n881), .A2(n880), .Z(n733) );
  XOR2D1BWP U1100 ( .A1(n944), .A2(n943), .Z(n945) );
  XOR2D1BWP U1101 ( .A1(n948), .A2(n949), .Z(n921) );
  XOR2D1BWP U1102 ( .A1(n869), .A2(n868), .Z(n874) );
  INVD3BWP U1480 ( .I(reset), .ZN(n1415) );
  INR2XD2BWP U1481 ( .A1(cu0_RegisterBlock_FF_io_data_out_1_), .B1(n1403), 
        .ZN(n740) );
  CKND1BWP U1482 ( .I(cu0_counterChain_io_data_0_out_1_), .ZN(n738) );
  IND2D1BWP U1483 ( .A1(n738), .B1(n1403), .ZN(n739) );
  CKND1BWP U1484 ( .I(cu0_RegisterBlock_FF_io_data_out_0_), .ZN(n741) );
  ND2D1BWP U1485 ( .A1(n1403), .A2(cu0_counterChain_io_data_0_out_0_), .ZN(
        n742) );
  AN2D1BWP U1486 ( .A1(n996), .A2(n743), .Z(cu0_RegisterBlock_FF_1_net3497) );
  ND2D1BWP U1487 ( .A1(n730), .A2(cu0_RegisterBlock_FF_io_data_out_6_), .ZN(
        n744) );
  FICIND1BWP U1488 ( .CIN(n744), .B(n730), .A(n730), .S(n745) );
  AN2D1BWP U1489 ( .A1(cu1_RegisterBlock_1_FF_1_io_data_out_7_), .A2(n1403), 
        .Z(n763) );
  ND2D1BWP U1490 ( .A1(n730), .A2(cu1_RegisterBlock_1_FF_io_data_out_5_), .ZN(
        n746) );
  IOA21D1BWP U1491 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_5_), 
        .B(n746), .ZN(n902) );
  CKND1BWP U1492 ( .I(cu1_RegisterBlock_io_passDataOut_1[5]), .ZN(n747) );
  OAI21D1BWP U1493 ( .A1(n730), .A2(n747), .B(n746), .ZN(n901) );
  IOA21D1BWP U1494 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_4_), 
        .B(n748), .ZN(n914) );
  CKND1BWP U1495 ( .I(cu1_RegisterBlock_io_passDataOut_1[4]), .ZN(n749) );
  OAI21D1BWP U1496 ( .A1(n730), .A2(n749), .B(n748), .ZN(n913) );
  ND2D1BWP U1497 ( .A1(n730), .A2(cu1_RegisterBlock_1_FF_io_data_out_3_), .ZN(
        n750) );
  IOA21D1BWP U1498 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_3_), 
        .B(n750), .ZN(n905) );
  CKND1BWP U1499 ( .I(cu1_RegisterBlock_io_passDataOut_1[3]), .ZN(n751) );
  OAI21D1BWP U1500 ( .A1(n730), .A2(n751), .B(n750), .ZN(n904) );
  IOA21D1BWP U1501 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_2_), 
        .B(n752), .ZN(n911) );
  CKND1BWP U1502 ( .I(cu1_RegisterBlock_io_passDataOut_1[2]), .ZN(n753) );
  OAI21D1BWP U1503 ( .A1(n730), .A2(n753), .B(n752), .ZN(n910) );
  ND2D1BWP U1504 ( .A1(n1403), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_1_), 
        .ZN(n754) );
  ND2D1BWP U1505 ( .A1(n724), .A2(n754), .ZN(n908) );
  ND2D1BWP U1506 ( .A1(n1403), .A2(cu1_RegisterBlock_io_passDataOut_1[1]), 
        .ZN(n755) );
  ND2D1BWP U1507 ( .A1(n724), .A2(n755), .ZN(n907) );
  INR2D2BWP U1508 ( .A1(cu1_RegisterBlock_1_FF_io_data_out_0_), .B1(n1403), 
        .ZN(n756) );
  CKND2BWP U1509 ( .I(n756), .ZN(n758) );
  ND2D1BWP U1510 ( .A1(n1403), .A2(cu1_RegisterBlock_io_passDataOut_1[0]), 
        .ZN(n757) );
  ND2D1BWP U1511 ( .A1(n758), .A2(n757), .ZN(n888) );
  ND2D1BWP U1512 ( .A1(n730), .A2(cu1_RegisterBlock_1_FF_io_data_out_6_), .ZN(
        n759) );
  AN2XD1BWP U1513 ( .A1(n766), .A2(n765), .Z(n760) );
  CKND4BWP U1514 ( .I(n764), .ZN(n887) );
  CKND6BWP U1515 ( .I(n887), .ZN(n1416) );
  XOR2D1BWP U1516 ( .A1(n766), .A2(n765), .Z(n767) );
  IND2D1BWP U1517 ( .A1(n1403), .B1(cu0_RegisterBlock_1_FF_io_data_out_0_), 
        .ZN(n771) );
  ND2D1BWP U1518 ( .A1(n1403), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_0_), 
        .ZN(n770) );
  ND2D1BWP U1519 ( .A1(n1403), .A2(cu1_counterChain_io_data_0_out_2_), .ZN(
        n772) );
  INR2XD1BWP U1520 ( .A1(cu1_RegisterBlock_FF_io_data_out_1_), .B1(n1403), 
        .ZN(n773) );
  CKND2BWP U1521 ( .I(n773), .ZN(n780) );
  ND2D1BWP U1522 ( .A1(n1403), .A2(cu1_counterChain_io_data_1_out_1_), .ZN(
        n774) );
  NR2D1BWP U1523 ( .A1(n932), .A2(n930), .ZN(n919) );
  CKND1BWP U1524 ( .I(cu1_RegisterBlock_FF_io_data_out_0_), .ZN(n775) );
  INR2D1BWP U1525 ( .A1(cu1_RegisterBlock_FF_io_data_out_3_), .B1(n1403), .ZN(
        n995) );
  NR2D1BWP U1526 ( .A1(n936), .A2(n942), .ZN(n918) );
  NR2D1BWP U1527 ( .A1(n936), .A2(n941), .ZN(n789) );
  INVD1BWP U1528 ( .I(cu1_counterChain_io_data_0_out_1_), .ZN(n779) );
  CKND2BWP U1529 ( .I(n839), .ZN(n931) );
  NR2D1BWP U1530 ( .A1(n931), .A2(n930), .ZN(n788) );
  NR2D1BWP U1531 ( .A1(n931), .A2(n941), .ZN(n916) );
  CKND1BWP U1532 ( .I(cu1_counterChain_io_data_1_out_0_), .ZN(n783) );
  NR2D1BWP U1533 ( .A1(n942), .A2(n937), .ZN(n915) );
  CKND1BWP U1534 ( .I(n924), .ZN(n787) );
  ND2D1BWP U1535 ( .A1(n786), .A2(n785), .ZN(n922) );
  ND2D1BWP U1536 ( .A1(n787), .A2(n922), .ZN(n793) );
  HA1D1BWP U1537 ( .A(n789), .B(n788), .CO(n917), .S(n791) );
  NR2D1BWP U1538 ( .A1(n932), .A2(n937), .ZN(n790) );
  OR2XD1BWP U1539 ( .A1(n791), .A2(n790), .Z(n819) );
  NR2D1BWP U1540 ( .A1(n931), .A2(n937), .ZN(n843) );
  NR2D1BWP U1541 ( .A1(n936), .A2(n930), .ZN(n842) );
  ND2D1BWP U1542 ( .A1(n843), .A2(n842), .ZN(n844) );
  CKND1BWP U1543 ( .I(n844), .ZN(n820) );
  ND2D1BWP U1544 ( .A1(n791), .A2(n790), .ZN(n818) );
  CKND1BWP U1545 ( .I(n818), .ZN(n792) );
  AOI21D1BWP U1546 ( .A1(n819), .A2(n820), .B(n792), .ZN(n923) );
  XOR2D1BWP U1547 ( .A1(n793), .A2(n923), .Z(cu1_IntFU_T7[3]) );
  ND2D1BWP U1548 ( .A1(cu1_IntFU_T7[3]), .A2(n726), .ZN(n796) );
  ND2D1BWP U1549 ( .A1(n794), .A2(n730), .ZN(n795) );
  AN2D1BWP U1550 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_7_), .A2(n726), 
        .Z(n814) );
  CKND1BWP U1551 ( .I(cu0_RegisterBlock_io_passDataOut_1[5]), .ZN(n798) );
  OAI21D1BWP U1552 ( .A1(n730), .A2(n798), .B(n797), .ZN(n891) );
  IOA21D2BWP U1553 ( .A1(n1403), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_4_), 
        .B(n799), .ZN(n899) );
  CKND1BWP U1554 ( .I(cu0_RegisterBlock_io_passDataOut_1[4]), .ZN(n800) );
  OAI21D1BWP U1555 ( .A1(n730), .A2(n800), .B(n799), .ZN(n898) );
  CKND1BWP U1556 ( .I(cu0_RegisterBlock_io_passDataOut_1[3]), .ZN(n802) );
  IOA21D1BWP U1557 ( .A1(n1403), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_2_), 
        .B(n803), .ZN(n896) );
  CKND1BWP U1558 ( .I(cu0_RegisterBlock_io_passDataOut_1[2]), .ZN(n804) );
  OAI21D1BWP U1559 ( .A1(n730), .A2(n804), .B(n803), .ZN(n895) );
  NR2D1BWP U1560 ( .A1(n806), .A2(n805), .ZN(n809) );
  CKND1BWP U1561 ( .I(n805), .ZN(n808) );
  CKND1BWP U1562 ( .I(n806), .ZN(n807) );
  AN2XD1BWP U1563 ( .A1(n811), .A2(n857), .Z(n812) );
  OAI22D1BWP U1564 ( .A1(n859), .A2(n812), .B1(n811), .B2(n857), .ZN(n813) );
  CKND6BWP U1565 ( .I(n732), .ZN(n1405) );
  FA1D1BWP U1566 ( .A(n817), .B(n816), .CI(n815), .CO(n794), .S(n822) );
  ND2D1BWP U1567 ( .A1(n819), .A2(n818), .ZN(n821) );
  XNR2D1BWP U1568 ( .A1(n821), .A2(n820), .ZN(n966) );
  FICOND1BWP U1569 ( .A(n825), .B(n826), .CI(n823), .CON(n882), .S(n831) );
  CKND2BWP U1570 ( .I(n825), .ZN(n861) );
  NR2D1BWP U1571 ( .A1(n846), .A2(n861), .ZN(n848) );
  NR2D1BWP U1572 ( .A1(n864), .A2(n860), .ZN(n847) );
  NR2D1BWP U1573 ( .A1(n862), .A2(n845), .ZN(n828) );
  OR2XD1BWP U1574 ( .A1(n829), .A2(n828), .Z(n855) );
  ND2D1BWP U1575 ( .A1(n829), .A2(n828), .ZN(n852) );
  ND2D1BWP U1576 ( .A1(n855), .A2(n852), .ZN(n830) );
  NR2D1BWP U1577 ( .A1(n864), .A2(n845), .ZN(n837) );
  NR2D1BWP U1578 ( .A1(n846), .A2(n860), .ZN(n836) );
  ND2D1BWP U1579 ( .A1(n837), .A2(n836), .ZN(n838) );
  CKND1BWP U1580 ( .I(n838), .ZN(n854) );
  XNR2D1BWP U1581 ( .A1(n830), .A2(n854), .ZN(n967) );
  NR2D1BWP U1582 ( .A1(n936), .A2(n937), .ZN(n963) );
  AN2D1BWP U1583 ( .A1(n963), .A2(n1403), .Z(n1407) );
  FICIND1BWP U1584 ( .CIN(n832), .B(n833), .A(n834), .CO(n823), .S(n835) );
  FICIND1BWP U1585 ( .CIN(n936), .B(n839), .A(n840), .CO(n815), .S(n841) );
  NR2D1BWP U1586 ( .A1(n846), .A2(n845), .ZN(n962) );
  AN2D1BWP U1587 ( .A1(n962), .A2(n1403), .Z(n1411) );
  NR2D1BWP U1588 ( .A1(n862), .A2(n860), .ZN(n872) );
  NR2D1BWP U1589 ( .A1(n846), .A2(n863), .ZN(n871) );
  HA1D1BWP U1590 ( .A(n848), .B(n847), .CO(n870), .S(n829) );
  CKND1BWP U1591 ( .I(n876), .ZN(n851) );
  ND2D1BWP U1592 ( .A1(n850), .A2(n849), .ZN(n875) );
  ND2D1BWP U1593 ( .A1(n851), .A2(n875), .ZN(n856) );
  CKND1BWP U1594 ( .I(n852), .ZN(n853) );
  AOI21D1BWP U1595 ( .A1(n855), .A2(n854), .B(n853), .ZN(n877) );
  XOR2D1BWP U1596 ( .A1(n856), .A2(n877), .Z(cu0_IntFU_T7[3]) );
  XNR2D1BWP U1597 ( .A1(n811), .A2(n857), .ZN(n858) );
  XOR2D2BWP U1598 ( .A1(n859), .A2(n858), .Z(n968) );
  CKND6BWP U1599 ( .I(n968), .ZN(n1404) );
  NR2D1BWP U1600 ( .A1(n863), .A2(n860), .ZN(n867) );
  NR2D1BWP U1601 ( .A1(n862), .A2(n861), .ZN(n866) );
  NR2D1BWP U1602 ( .A1(n864), .A2(n863), .ZN(n865) );
  FA1D1BWP U1603 ( .A(n867), .B(n866), .CI(n865), .S(n868) );
  FA1D1BWP U1604 ( .A(n872), .B(n871), .CI(n870), .CO(n873), .S(n850) );
  ND2D1BWP U1605 ( .A1(n874), .A2(n873), .ZN(n954) );
  CKND1BWP U1606 ( .I(n954), .ZN(n881) );
  OR2XD1BWP U1607 ( .A1(n874), .A2(n873), .Z(n955) );
  OAI21D1BWP U1608 ( .A1(n877), .A2(n876), .B(n875), .ZN(n956) );
  CKND1BWP U1609 ( .I(n956), .ZN(n878) );
  ND2D1BWP U1610 ( .A1(n733), .A2(n1406), .ZN(n969) );
  CKND1BWP U1611 ( .I(n969), .ZN(cu0_RegisterBlock_FF_3_net3500) );
  ND2D1BWP U1612 ( .A1(cu0_IntFU_T7[3]), .A2(n1403), .ZN(n886) );
  FICIND1BWP U1613 ( .CIN(n882), .B(n883), .A(n883), .CO(n997), .S(n884) );
  ND2D1BWP U1614 ( .A1(n884), .A2(n730), .ZN(n885) );
  CKND1BWP U1615 ( .I(n996), .ZN(cu1_RegisterBlock_1_FF_1_net3491) );
  FICIND2BWP U1616 ( .CIN(n890), .B(n891), .A(n892), .CO(n859), .S(
        cu0_IntFU_1_m_T3[5]) );
  FICOND2BWP U1617 ( .A(n896), .B(n895), .CI(n894), .CON(n893), .S(
        cu0_IntFU_1_m_T3[2]) );
  FICOND2BWP U1618 ( .A(n899), .B(n898), .CI(n897), .CON(n890), .S(
        cu0_IntFU_1_m_T3[4]) );
  FICIND2BWP U1619 ( .CIN(n900), .B(n901), .A(n902), .CO(n768), .S(
        cu1_IntFU_1_m_T3[5]) );
  FICIND2BWP U1620 ( .CIN(n903), .B(n904), .A(n905), .CO(n912), .S(
        cu1_IntFU_1_m_T3[3]) );
  FICIND2BWP U1621 ( .CIN(n906), .B(n907), .A(n908), .CO(n909), .S(
        cu1_IntFU_1_m_T3[1]) );
  FICOND2BWP U1622 ( .A(n911), .B(n910), .CI(n909), .CON(n903), .S(
        cu1_IntFU_1_m_T3[2]) );
  FICOND2BWP U1623 ( .A(n914), .B(n913), .CI(n912), .CON(n900), .S(
        cu1_IntFU_1_m_T3[4]) );
  HA1D1BWP U1624 ( .A(n916), .B(n915), .CO(n949), .S(n785) );
  NR2D1BWP U1625 ( .A1(n942), .A2(n930), .ZN(n928) );
  NR2D1BWP U1626 ( .A1(n932), .A2(n941), .ZN(n927) );
  NR2D1BWP U1627 ( .A1(n931), .A2(n942), .ZN(n926) );
  ND2D1BWP U1628 ( .A1(n921), .A2(n920), .ZN(n951) );
  ND2D1BWP U1629 ( .A1(n952), .A2(n951), .ZN(n925) );
  OAI21D1BWP U1630 ( .A1(n924), .A2(n923), .B(n922), .ZN(n953) );
  XNR2D1BWP U1631 ( .A1(n925), .A2(n953), .ZN(cu1_IntFU_T7[4]) );
  FA1D1BWP U1632 ( .A(n928), .B(n927), .CI(n926), .CO(n947), .S(n948) );
  NR2D1BWP U1633 ( .A1(n938), .A2(n930), .ZN(n935) );
  NR2D1BWP U1634 ( .A1(n931), .A2(n938), .ZN(n934) );
  NR2D1BWP U1635 ( .A1(n932), .A2(n942), .ZN(n933) );
  NR2D1BWP U1636 ( .A1(n936), .A2(n938), .ZN(n940) );
  NR2D1BWP U1637 ( .A1(n938), .A2(n937), .ZN(n939) );
  NR2D1BWP U1638 ( .A1(n942), .A2(n941), .ZN(n943) );
  ND2D1BWP U1639 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNR2D1BWP U1640 ( .A1(n957), .A2(n956), .ZN(cu0_IntFU_T7[4]) );
  AN2XD1BWP U1641 ( .A1(io_command), .A2(n1415), .Z(controlBox_N6) );
  XNR2D1BWP U1642 ( .A1(cu0_counterChain_io_data_1_out_0_), .A2(
        cu0_counterChain_io_data_1_out_1_), .ZN(n958) );
  NR2D1BWP U1643 ( .A1(n958), .A2(n1020), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net3512) );
  XNR2D1BWP U1644 ( .A1(cu1_counterChain_io_data_1_out_0_), .A2(
        cu1_counterChain_io_data_1_out_1_), .ZN(n959) );
  NR2D1BWP U1645 ( .A1(n959), .A2(n1024), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net3512) );
  XNR2D1BWP U1646 ( .A1(cu0_counterChain_io_data_0_out_0_), .A2(
        cu0_counterChain_io_data_0_out_1_), .ZN(n960) );
  NR2D1BWP U1647 ( .A1(n960), .A2(n1018), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net3512) );
  XNR2D1BWP U1648 ( .A1(cu1_counterChain_io_data_0_out_0_), .A2(
        cu1_counterChain_io_data_0_out_1_), .ZN(n961) );
  NR2D1BWP U1649 ( .A1(n961), .A2(n1022), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net3512) );
  AO22D1BWP U1650 ( .A1(n962), .A2(n1406), .B1(n996), .B2(
        cu0_counterChain_io_data_1_out_0_), .Z(cu0_RegisterBlock_FF_3_net3515)
         );
  AO22D1BWP U1651 ( .A1(n963), .A2(n1406), .B1(n996), .B2(
        cu1_counterChain_io_data_1_out_0_), .Z(cu1_RegisterBlock_FF_3_net3515)
         );
  AO22D1BWP U1652 ( .A1(n964), .A2(n1406), .B1(n996), .B2(
        cu0_counterChain_io_data_1_out_1_), .Z(cu0_RegisterBlock_FF_3_net3512)
         );
  AO22D1BWP U1653 ( .A1(n965), .A2(n1406), .B1(n996), .B2(
        cu1_counterChain_io_data_1_out_1_), .Z(cu1_RegisterBlock_FF_3_net3512)
         );
  AO22D1BWP U1654 ( .A1(n966), .A2(n1406), .B1(n996), .B2(
        cu1_counterChain_io_data_1_out_2_), .Z(cu1_RegisterBlock_FF_3_net3509)
         );
  AO22D1BWP U1655 ( .A1(n967), .A2(n1406), .B1(n996), .B2(
        cu0_counterChain_io_data_1_out_2_), .Z(cu0_RegisterBlock_FF_3_net3509)
         );
  NR2D1BWP U1656 ( .A1(n968), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_1_net3497) );
  IOA21D1BWP U1657 ( .A1(n970), .A2(n996), .B(n969), .ZN(
        cu0_RegisterBlock_FF_1_net3500) );
  CKND1BWP U1658 ( .I(n1410), .ZN(n971) );
  NR2D1BWP U1659 ( .A1(reset), .A2(n971), .ZN(cu1_RegisterBlock_FF_1_net3506)
         );
  CKND1BWP U1660 ( .I(n1411), .ZN(n973) );
  NR2D1BWP U1661 ( .A1(n974), .A2(n979), .ZN(cu0_mem0_N23) );
  INR2D1BWP U1662 ( .A1(n1411), .B1(n1412), .ZN(n972) );
  INVD1BWP U1663 ( .I(n972), .ZN(n977) );
  NR2D1BWP U1664 ( .A1(n974), .A2(n977), .ZN(cu0_mem0_N24) );
  ND2D1BWP U1665 ( .A1(n1412), .A2(n973), .ZN(n980) );
  NR2D1BWP U1666 ( .A1(n974), .A2(n980), .ZN(cu0_mem0_N25) );
  INVD1BWP U1667 ( .I(n975), .ZN(n976) );
  ND2D1BWP U1668 ( .A1(n1412), .A2(n1411), .ZN(n981) );
  NR2D1BWP U1669 ( .A1(n976), .A2(n981), .ZN(cu0_mem0_N22) );
  NR2D1BWP U1670 ( .A1(n977), .A2(n976), .ZN(cu0_mem0_N20) );
  NR2D1BWP U1671 ( .A1(n979), .A2(n976), .ZN(cu0_mem0_N19) );
  NR2D1BWP U1672 ( .A1(n980), .A2(n976), .ZN(cu0_mem0_N21) );
  NR2D1BWP U1673 ( .A1(n978), .A2(n979), .ZN(cu0_mem0_N15) );
  NR2D1BWP U1674 ( .A1(n978), .A2(n977), .ZN(cu0_mem0_N16) );
  NR2D1BWP U1675 ( .A1(n978), .A2(n980), .ZN(cu0_mem0_N17) );
  NR2D1BWP U1676 ( .A1(n978), .A2(n981), .ZN(cu0_mem0_N18) );
  ND2D1BWP U1677 ( .A1(n1414), .A2(n1413), .ZN(n982) );
  NR2D1BWP U1678 ( .A1(n982), .A2(n979), .ZN(cu0_mem0_N27) );
  NR2D1BWP U1679 ( .A1(n982), .A2(n980), .ZN(cu0_mem0_N29) );
  NR2D1BWP U1680 ( .A1(n982), .A2(n981), .ZN(cu0_mem0_N30) );
  NR2D1BWP U1681 ( .A1(n732), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_1_net3494) );
  INR2XD1BWP U1682 ( .A1(n1409), .B1(n1410), .ZN(n983) );
  ND2D1BWP U1683 ( .A1(n1408), .A2(n1407), .ZN(n988) );
  NR2D1BWP U1684 ( .A1(n985), .A2(n988), .ZN(cu1_mem1_N22) );
  CKND1BWP U1685 ( .I(n1407), .ZN(n984) );
  NR2D1BWP U1686 ( .A1(n993), .A2(n985), .ZN(cu1_mem1_N19) );
  NR2D1BWP U1687 ( .A1(n990), .A2(n985), .ZN(cu1_mem1_N20) );
  ND2D1BWP U1688 ( .A1(n1408), .A2(n984), .ZN(n992) );
  NR2D1BWP U1689 ( .A1(n992), .A2(n985), .ZN(cu1_mem1_N21) );
  CKND1BWP U1690 ( .I(n1409), .ZN(n989) );
  NR2D1BWP U1691 ( .A1(n987), .A2(n993), .ZN(cu1_mem1_N15) );
  NR2D1BWP U1692 ( .A1(n987), .A2(n990), .ZN(cu1_mem1_N16) );
  NR2D1BWP U1693 ( .A1(n987), .A2(n992), .ZN(cu1_mem1_N17) );
  NR2D1BWP U1694 ( .A1(n987), .A2(n988), .ZN(cu1_mem1_N18) );
  ND2D1BWP U1696 ( .A1(n1410), .A2(n1409), .ZN(n994) );
  NR2D1BWP U1697 ( .A1(n994), .A2(n988), .ZN(cu1_mem1_N30) );
  ND2D1BWP U1698 ( .A1(n1410), .A2(n989), .ZN(n991) );
  NR2D1BWP U1699 ( .A1(n991), .A2(n990), .ZN(cu1_mem1_N24) );
  NR2D1BWP U1700 ( .A1(n991), .A2(n993), .ZN(cu1_mem1_N23) );
  NR2D1BWP U1701 ( .A1(n991), .A2(n992), .ZN(cu1_mem1_N25) );
  NR2D1BWP U1702 ( .A1(n994), .A2(n992), .ZN(cu1_mem1_N29) );
  NR2D1BWP U1703 ( .A1(n994), .A2(n993), .ZN(cu1_mem1_N27) );
  IND2D1BWP U1705 ( .A1(io_config_enable), .B1(n1415), .ZN(
        cu0_controlBlock_incXbar_net3599) );
  NR2D1BWP U1706 ( .A1(reset), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3581) );
  INR2D1BWP U1707 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__net3581), .B1(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n998) );
  AO31D1BWP U1708 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), 
        .A2(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n1415), .B(
        n998), .Z(cu1_controlBlock_UpDownCtr_1_reg__net3578) );
  NR2D1BWP U1709 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n1000) );
  CKND1BWP U1710 ( .I(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n999) );
  ND2D1BWP U1711 ( .A1(n998), .A2(n999), .ZN(n1002) );
  OAI31D1BWP U1712 ( .A1(reset), .A2(n1000), .A3(n999), .B(n1002), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3575) );
  OAI31D1BWP U1713 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n1001) );
  OAI22D1BWP U1714 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n1002), .B1(reset), .B2(n1001), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net3572) );
  NR2D1BWP U1715 ( .A1(reset), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3581) );
  INR2D1BWP U1716 ( .A1(cu0_controlBlock_UpDownCtr_reg__net3581), .B1(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n1003) );
  AO31D1BWP U1717 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n1415), .B(n1003), 
        .Z(cu0_controlBlock_UpDownCtr_reg__net3578) );
  NR2D1BWP U1718 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n1005) );
  CKND1BWP U1719 ( .I(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(
        n1004) );
  ND2D1BWP U1720 ( .A1(n1003), .A2(n1004), .ZN(n1007) );
  OAI31D1BWP U1721 ( .A1(reset), .A2(n1005), .A3(n1004), .B(n1007), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3575) );
  OAI31D1BWP U1722 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n1006) );
  OAI22D1BWP U1723 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n1007), .B1(reset), .B2(n1006), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net3572) );
  NR2D1BWP U1724 ( .A1(reset), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3581) );
  INR2D1BWP U1725 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__net3581), .B1(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n1008) );
  AO31D1BWP U1726 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), 
        .A2(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n1415), .B(
        n1008), .Z(cu0_controlBlock_UpDownCtr_1_reg__net3578) );
  NR2D1BWP U1727 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n1010) );
  CKND1BWP U1728 ( .I(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n1009) );
  ND2D1BWP U1729 ( .A1(n1008), .A2(n1009), .ZN(n1012) );
  OAI31D1BWP U1730 ( .A1(reset), .A2(n1010), .A3(n1009), .B(n1012), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3575) );
  OAI31D1BWP U1731 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n1011) );
  OAI22D1BWP U1732 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n1012), .B1(reset), .B2(n1011), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net3572) );
  NR2D1BWP U1733 ( .A1(reset), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3581) );
  INR2D1BWP U1734 ( .A1(cu1_controlBlock_UpDownCtr_reg__net3581), .B1(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n1013) );
  AO31D1BWP U1735 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n1415), .B(n1013), 
        .Z(cu1_controlBlock_UpDownCtr_reg__net3578) );
  NR2D1BWP U1736 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n1015) );
  CKND1BWP U1737 ( .I(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(
        n1014) );
  ND2D1BWP U1738 ( .A1(n1013), .A2(n1014), .ZN(n1017) );
  OAI31D1BWP U1739 ( .A1(reset), .A2(n1015), .A3(n1014), .B(n1017), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3575) );
  OAI31D1BWP U1740 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n1016) );
  OAI22D1BWP U1741 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n1017), .B1(reset), .B2(n1016), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net3572) );
  NR2D1BWP U1742 ( .A1(n1018), .A2(cu0_counterChain_io_data_0_out_0_), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net3515) );
  CKND2D1BWP U1743 ( .A1(cu0_counterChain_io_data_0_out_0_), .A2(
        cu0_counterChain_io_data_0_out_1_), .ZN(n1019) );
  NR2D1BWP U1744 ( .A1(n1019), .A2(n1018), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net3509) );
  NR2D1BWP U1745 ( .A1(n1020), .A2(cu0_counterChain_io_data_1_out_0_), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net3515) );
  CKND2D1BWP U1746 ( .A1(cu0_counterChain_io_data_1_out_0_), .A2(
        cu0_counterChain_io_data_1_out_1_), .ZN(n1021) );
  NR2D1BWP U1747 ( .A1(n1021), .A2(n1020), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net3509) );
  NR2D1BWP U1748 ( .A1(n1022), .A2(cu1_counterChain_io_data_0_out_0_), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net3515) );
  CKND2D1BWP U1749 ( .A1(cu1_counterChain_io_data_0_out_0_), .A2(
        cu1_counterChain_io_data_0_out_1_), .ZN(n1023) );
  NR2D1BWP U1750 ( .A1(n1023), .A2(n1022), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net3509) );
  NR2D1BWP U1751 ( .A1(n1024), .A2(cu1_counterChain_io_data_1_out_0_), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net3515) );
  CKND2D1BWP U1752 ( .A1(cu1_counterChain_io_data_1_out_0_), .A2(
        cu1_counterChain_io_data_1_out_1_), .ZN(n1025) );
  NR2D1BWP U1753 ( .A1(n1025), .A2(n1024), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net3509) );
endmodule

