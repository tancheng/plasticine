
module SRAM ( clk, io_raddr, io_wen, io_waddr, io_wdata, io_rdata );
  input [3:0] io_raddr;
  input [3:0] io_waddr;
  input [7:0] io_wdata;
  output [7:0] io_rdata;
  input clk, io_wen;


endmodule


module SNPS_CLOCK_GATE_HIGH_FF_1_4_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_FF_1_4_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CKLNQD1BWP latch ( .CP(CLK), .E(EN), .TE(TE), .Q(ENCLK) );
endmodule


module Plasticine ( clk, reset, io_config_enable, io_command, io_status );
  input clk, reset, io_config_enable, io_command;
  output io_status;
  wire   controlBox_N6, controlBox_commandReg,
         cu1_counterChain_io_data_0_out_0_, cu1_counterChain_io_data_0_out_1_,
         cu1_counterChain_io_data_0_out_2_, cu1_counterChain_io_data_1_out_0_,
         cu1_counterChain_io_data_1_out_1_, cu1_counterChain_io_data_1_out_2_,
         cu1_mem1_io_rdata_0_, cu1_mem1_io_rdata_1_, cu1_mem1_io_rdata_2_,
         cu1_mem1_io_rdata_3_, cu1_mem1_io_rdata_4_, cu1_mem1_io_rdata_5_,
         cu1_mem1_io_rdata_6_, cu1_mem1_io_rdata_7_, cu1_mem0_io_rdata_0_,
         cu1_mem0_io_rdata_1_, cu1_mem0_io_rdata_2_, cu1_mem0_io_rdata_3_,
         cu1_mem0_io_rdata_4_, cu1_mem0_io_rdata_5_, cu1_mem0_io_rdata_6_,
         cu1_mem0_io_rdata_7_, cu0_counterChain_io_data_0_out_0_,
         cu0_counterChain_io_data_0_out_1_, cu0_counterChain_io_data_0_out_2_,
         cu0_counterChain_io_data_1_out_0_, cu0_counterChain_io_data_1_out_1_,
         cu0_counterChain_io_data_1_out_2_, cu0_mem1_io_rdata_0_,
         cu0_mem1_io_rdata_1_, cu0_mem1_io_rdata_2_, cu0_mem1_io_rdata_3_,
         cu0_mem1_io_rdata_4_, cu0_mem1_io_rdata_5_, cu0_mem1_io_rdata_6_,
         cu0_mem1_io_rdata_7_, cu0_mem0_io_rdata_0_, cu0_mem0_io_rdata_1_,
         cu0_mem0_io_rdata_2_, cu0_mem0_io_rdata_3_, cu0_mem0_io_rdata_4_,
         cu0_mem0_io_rdata_5_, cu0_mem0_io_rdata_6_, cu0_mem0_io_rdata_7_,
         cu0_T21_0_, controlBox_pulser_N3,
         cu1_RegisterBlock_1_FF_1_io_data_out_0_,
         cu1_RegisterBlock_1_FF_1_io_data_out_1_,
         cu1_RegisterBlock_1_FF_1_io_data_out_2_,
         cu1_RegisterBlock_1_FF_1_io_data_out_3_,
         cu1_RegisterBlock_1_FF_1_io_data_out_4_,
         cu1_RegisterBlock_1_FF_1_io_data_out_5_,
         cu1_RegisterBlock_1_FF_1_io_data_out_6_,
         cu1_RegisterBlock_1_FF_1_io_data_out_7_,
         cu1_RegisterBlock_1_FF_io_data_out_0_,
         cu1_RegisterBlock_1_FF_io_data_out_1_,
         cu1_RegisterBlock_1_FF_io_data_out_2_,
         cu1_RegisterBlock_1_FF_io_data_out_3_,
         cu1_RegisterBlock_1_FF_io_data_out_4_,
         cu1_RegisterBlock_1_FF_io_data_out_5_,
         cu1_RegisterBlock_1_FF_io_data_out_6_,
         cu1_RegisterBlock_FF_io_data_out_0_,
         cu1_RegisterBlock_FF_io_data_out_1_,
         cu1_RegisterBlock_FF_io_data_out_2_,
         cu1_RegisterBlock_FF_io_data_out_3_,
         cu1_RegisterBlock_FF_io_data_out_4_,
         cu1_RegisterBlock_FF_io_data_out_5_,
         cu1_RegisterBlock_FF_io_data_out_6_,
         cu0_RegisterBlock_FF_io_data_out_0_,
         cu0_RegisterBlock_FF_io_data_out_1_,
         cu0_RegisterBlock_FF_io_data_out_2_,
         cu0_RegisterBlock_FF_io_data_out_3_,
         cu0_RegisterBlock_FF_io_data_out_4_,
         cu0_RegisterBlock_FF_io_data_out_5_,
         cu0_RegisterBlock_FF_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_0_,
         cu0_RegisterBlock_1_FF_1_io_data_out_1_,
         cu0_RegisterBlock_1_FF_1_io_data_out_2_,
         cu0_RegisterBlock_1_FF_1_io_data_out_3_,
         cu0_RegisterBlock_1_FF_1_io_data_out_4_,
         cu0_RegisterBlock_1_FF_1_io_data_out_5_,
         cu0_RegisterBlock_1_FF_1_io_data_out_6_,
         cu0_RegisterBlock_1_FF_1_io_data_out_7_,
         cu0_RegisterBlock_1_FF_io_data_out_0_,
         cu0_RegisterBlock_1_FF_io_data_out_1_,
         cu0_RegisterBlock_1_FF_io_data_out_2_,
         cu0_RegisterBlock_1_FF_io_data_out_3_,
         cu0_RegisterBlock_1_FF_io_data_out_4_,
         cu0_RegisterBlock_1_FF_io_data_out_5_,
         cu0_RegisterBlock_1_FF_io_data_out_6_,
         cu1_RegisterBlock_1_FF_5_net4412, cu1_RegisterBlock_1_FF_5_net4409,
         cu1_RegisterBlock_1_FF_5_net4406, cu1_RegisterBlock_1_FF_5_net4403,
         cu1_RegisterBlock_1_FF_5_net4400, cu1_RegisterBlock_1_FF_5_net4397,
         cu1_RegisterBlock_1_FF_5_net4394,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu1_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_incXbar_net4499, cu0_controlBlock_incXbar_net4496,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_reg__io_data_out_3_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_,
         cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_,
         cu0_RegisterBlock_FF_1_net4412, cu0_RegisterBlock_FF_1_net4409,
         cu0_RegisterBlock_FF_1_net4406, cu0_RegisterBlock_FF_1_net4403,
         cu0_RegisterBlock_FF_1_net4400, cu0_RegisterBlock_FF_1_net4397,
         cu0_RegisterBlock_FF_2_net4412, cu0_RegisterBlock_FF_2_net4409,
         cu0_RegisterBlock_FF_2_net4406, cu0_RegisterBlock_FF_3_net4412,
         cu0_RegisterBlock_FF_3_net4409, cu0_RegisterBlock_FF_3_net4406,
         cu0_RegisterBlock_FF_3_net4403, cu0_RegisterBlock_FF_3_net4400,
         cu0_RegisterBlock_FF_3_net4397, cu0_RegisterBlock_FF_4_net4412,
         cu0_RegisterBlock_FF_4_net4409, cu0_RegisterBlock_FF_4_net4406,
         cu0_RegisterBlock_FF_4_net4403, cu0_RegisterBlock_FF_4_net4400,
         cu0_RegisterBlock_FF_4_net4397, cu0_RegisterBlock_FF_4_net4394,
         cu0_RegisterBlock_FF_4_net4391, cu0_RegisterBlock_FF_5_net4412,
         cu0_RegisterBlock_FF_5_net4409, cu0_RegisterBlock_FF_5_net4406,
         cu0_RegisterBlock_FF_5_net4403, cu0_RegisterBlock_FF_5_net4400,
         cu0_RegisterBlock_FF_5_net4397, cu0_RegisterBlock_FF_5_net4394,
         cu0_RegisterBlock_FF_5_net4391, cu0_RegisterBlock_1_FF_1_net4412,
         cu0_RegisterBlock_1_FF_1_net4409, cu0_RegisterBlock_1_FF_1_net4406,
         cu0_RegisterBlock_1_FF_1_net4403, cu0_RegisterBlock_1_FF_1_net4400,
         cu0_RegisterBlock_1_FF_1_net4397, cu0_RegisterBlock_1_FF_1_net4394,
         cu0_RegisterBlock_1_FF_1_net4391, cu0_RegisterBlock_1_FF_2_net4412,
         cu0_RegisterBlock_1_FF_2_net4409, cu0_RegisterBlock_1_FF_2_net4406,
         cu0_RegisterBlock_1_FF_3_net4412, cu0_RegisterBlock_1_FF_3_net4409,
         cu0_RegisterBlock_1_FF_3_net4406, cu0_RegisterBlock_1_FF_3_net4403,
         cu0_RegisterBlock_1_FF_3_net4400, cu0_RegisterBlock_1_FF_3_net4397,
         cu0_RegisterBlock_1_FF_4_net4412, cu0_RegisterBlock_1_FF_4_net4409,
         cu0_RegisterBlock_1_FF_4_net4406, cu0_RegisterBlock_1_FF_4_net4403,
         cu0_RegisterBlock_1_FF_4_net4400, cu0_RegisterBlock_1_FF_4_net4397,
         cu0_RegisterBlock_1_FF_4_net4394, cu0_RegisterBlock_1_FF_4_net4391,
         cu0_RegisterBlock_1_FF_5_net4412, cu0_RegisterBlock_1_FF_5_net4409,
         cu0_RegisterBlock_1_FF_5_net4406, cu0_RegisterBlock_1_FF_5_net4403,
         cu0_RegisterBlock_1_FF_5_net4400, cu0_RegisterBlock_1_FF_5_net4397,
         cu0_RegisterBlock_1_FF_5_net4394, cu0_RegisterBlock_1_FF_5_net4391,
         cu1_counterChain_CounterRC_config__stride_0_,
         cu1_RegisterBlock_FF_1_net4412, cu1_RegisterBlock_FF_1_net4409,
         cu1_RegisterBlock_FF_1_net4406, cu1_RegisterBlock_FF_1_net4403,
         cu1_RegisterBlock_FF_1_net4400, cu1_RegisterBlock_FF_1_net4397,
         cu1_RegisterBlock_FF_1_net4394, cu1_RegisterBlock_FF_2_net4412,
         cu1_RegisterBlock_FF_2_net4409, cu1_RegisterBlock_FF_3_net4412,
         cu1_RegisterBlock_FF_3_net4409, cu1_RegisterBlock_FF_3_net4406,
         cu1_RegisterBlock_FF_3_net4403, cu1_RegisterBlock_FF_3_net4400,
         cu1_RegisterBlock_FF_3_net4397, cu1_RegisterBlock_FF_4_net4412,
         cu1_RegisterBlock_FF_4_net4409, cu1_RegisterBlock_FF_4_net4406,
         cu1_RegisterBlock_FF_4_net4403, cu1_RegisterBlock_FF_4_net4400,
         cu1_RegisterBlock_FF_4_net4397, cu1_RegisterBlock_FF_4_net4394,
         cu1_RegisterBlock_FF_4_net4391, cu1_RegisterBlock_FF_5_net4412,
         cu1_RegisterBlock_FF_5_net4409, cu1_RegisterBlock_FF_5_net4406,
         cu1_RegisterBlock_FF_5_net4403, cu1_RegisterBlock_FF_5_net4400,
         cu1_RegisterBlock_FF_5_net4397, cu1_RegisterBlock_FF_5_net4394,
         cu1_RegisterBlock_FF_5_net4391, cu1_RegisterBlock_1_FF_1_net4415,
         cu1_RegisterBlock_1_FF_1_net4412, cu1_RegisterBlock_1_FF_1_net4409,
         cu1_RegisterBlock_1_FF_1_net4406, cu1_RegisterBlock_1_FF_1_net4403,
         cu1_RegisterBlock_1_FF_1_net4400, cu1_RegisterBlock_1_FF_1_net4397,
         cu1_RegisterBlock_1_FF_1_net4394, cu1_RegisterBlock_1_FF_1_net4391,
         cu1_RegisterBlock_1_FF_1_net4388, cu1_RegisterBlock_1_FF_2_net4412,
         cu1_RegisterBlock_1_FF_2_net4409, cu1_RegisterBlock_1_FF_2_net4406,
         cu1_RegisterBlock_1_FF_3_net4412, cu1_RegisterBlock_1_FF_3_net4409,
         cu1_RegisterBlock_1_FF_3_net4406, cu1_RegisterBlock_1_FF_3_net4403,
         cu1_RegisterBlock_1_FF_3_net4400, cu1_RegisterBlock_1_FF_3_net4397,
         cu1_RegisterBlock_1_FF_4_net4412, cu1_RegisterBlock_1_FF_4_net4409,
         cu1_RegisterBlock_1_FF_4_net4406, cu1_RegisterBlock_1_FF_4_net4403,
         cu1_RegisterBlock_1_FF_4_net4400, cu1_RegisterBlock_1_FF_4_net4397,
         cu1_RegisterBlock_1_FF_4_net4394, cu1_RegisterBlock_1_FF_4_net4391,
         cu1_controlBlock_UpDownCtr_1_reg__net4478,
         cu1_controlBlock_UpDownCtr_1_reg__net4475,
         cu1_controlBlock_UpDownCtr_1_reg__net4472,
         cu1_controlBlock_UpDownCtr_1_reg__net4469,
         cu0_controlBlock_UpDownCtr_reg__net4478,
         cu0_controlBlock_UpDownCtr_reg__net4475,
         cu0_controlBlock_UpDownCtr_reg__net4472,
         cu0_controlBlock_UpDownCtr_reg__net4469,
         cu0_controlBlock_UpDownCtr_1_reg__net4478,
         cu0_controlBlock_UpDownCtr_1_reg__net4475,
         cu0_controlBlock_UpDownCtr_1_reg__net4472,
         cu0_controlBlock_UpDownCtr_1_reg__net4469,
         cu1_controlBlock_UpDownCtr_reg__net4478,
         cu1_controlBlock_UpDownCtr_reg__net4475,
         cu1_controlBlock_UpDownCtr_reg__net4472,
         cu1_controlBlock_UpDownCtr_reg__net4469,
         cu0_counterChain_CounterRC_counter_reg__net4412,
         cu0_counterChain_CounterRC_counter_reg__net4409,
         cu0_counterChain_CounterRC_counter_reg__net4406,
         cu0_counterChain_CounterRC_1_counter_reg__net4412,
         cu0_counterChain_CounterRC_1_counter_reg__net4409,
         cu0_counterChain_CounterRC_1_counter_reg__net4406,
         cu1_counterChain_CounterRC_counter_reg__net4412,
         cu1_counterChain_CounterRC_counter_reg__net4409,
         cu1_counterChain_CounterRC_counter_reg__net4406,
         cu1_counterChain_CounterRC_1_counter_reg__net4415,
         cu1_counterChain_CounterRC_1_counter_reg__net4412,
         cu1_counterChain_CounterRC_1_counter_reg__net4409,
         cu1_counterChain_CounterRC_1_counter_reg__net4406, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333;
  wire   [2:0] cu1_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu1_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu1_RegisterBlock_io_passDataOut_2;
  wire   [7:0] cu1_RegisterBlock_io_passDataOut_3;
  wire   [3:0] cu1_mem0raMux_io_out_0;
  wire   [2:0] cu0_RegisterBlock_io_passDataOut_0;
  wire   [5:0] cu0_RegisterBlock_io_passDataOut_1;
  wire   [7:0] cu0_RegisterBlock_io_passDataOut_2;
  wire   [7:0] cu0_RegisterBlock_io_passDataOut_3;
  wire   [3:0] cu0_mem1raMux_io_out_0;
  wire   [7:0] cu1_IntFU_1_m_T3;
  wire   [7:0] cu0_IntFU_1_m_T3;
  assign io_status = 1'b0;

  SRAM cu1_mem1 ( .clk(clk), .io_raddr(cu1_mem0raMux_io_out_0), .io_wen(1'b1), 
        .io_waddr(cu1_mem0raMux_io_out_0), .io_wdata(cu1_IntFU_1_m_T3), 
        .io_rdata({cu1_mem1_io_rdata_7_, cu1_mem1_io_rdata_6_, 
        cu1_mem1_io_rdata_5_, cu1_mem1_io_rdata_4_, cu1_mem1_io_rdata_3_, 
        cu1_mem1_io_rdata_2_, cu1_mem1_io_rdata_1_, cu1_mem1_io_rdata_0_}) );
  SRAM cu1_mem0 ( .clk(clk), .io_raddr(cu1_mem0raMux_io_out_0), .io_wen(1'b1), 
        .io_waddr(cu1_mem0raMux_io_out_0), .io_wdata(cu1_IntFU_1_m_T3), 
        .io_rdata({cu1_mem0_io_rdata_7_, cu1_mem0_io_rdata_6_, 
        cu1_mem0_io_rdata_5_, cu1_mem0_io_rdata_4_, cu1_mem0_io_rdata_3_, 
        cu1_mem0_io_rdata_2_, cu1_mem0_io_rdata_1_, cu1_mem0_io_rdata_0_}) );
  SRAM cu0_mem1 ( .clk(clk), .io_raddr(cu0_mem1raMux_io_out_0), .io_wen(1'b1), 
        .io_waddr(cu0_mem1raMux_io_out_0), .io_wdata(cu0_IntFU_1_m_T3), 
        .io_rdata({cu0_mem1_io_rdata_7_, cu0_mem1_io_rdata_6_, 
        cu0_mem1_io_rdata_5_, cu0_mem1_io_rdata_4_, cu0_mem1_io_rdata_3_, 
        cu0_mem1_io_rdata_2_, cu0_mem1_io_rdata_1_, cu0_mem1_io_rdata_0_}) );
  SRAM cu0_mem0 ( .clk(clk), .io_raddr(cu0_mem1raMux_io_out_0), .io_wen(1'b1), 
        .io_waddr(cu0_mem1raMux_io_out_0), .io_wdata(cu0_IntFU_1_m_T3), 
        .io_rdata({cu0_mem0_io_rdata_7_, cu0_mem0_io_rdata_6_, 
        cu0_mem0_io_rdata_5_, cu0_mem0_io_rdata_4_, cu0_mem0_io_rdata_3_, 
        cu0_mem0_io_rdata_2_, cu0_mem0_io_rdata_1_, cu0_mem0_io_rdata_0_}) );
  SNPS_CLOCK_GATE_HIGH_Crossbar_1_0_1 cu0_controlBlock_incXbar_clk_gate_config__outSelect_3_reg ( 
        .CLK(clk), .EN(cu0_controlBlock_incXbar_net4496), .ENCLK(
        cu0_controlBlock_incXbar_net4499), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_8 cu1_RegisterBlock_1_FF_1_clk_gate_ff_reg ( 
        .CLK(clk), .EN(cu1_RegisterBlock_1_FF_1_net4388), .ENCLK(
        cu1_RegisterBlock_1_FF_1_net4415), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_FF_1_4_1 cu1_counterChain_CounterRC_1_counter_reg__clk_gate_ff_reg ( 
        .CLK(clk), .EN(reset), .ENCLK(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .TE(1'b0) );
  DFQD4BWP cu0_config__pipeStage_1_opB_value_reg_0_ ( .D(n332), .CP(
        cu0_controlBlock_incXbar_net4499), .Q(cu0_T21_0_) );
  DFQD4BWP controlBox_pulser_commandReg_reg ( .D(controlBox_pulser_N3), .CP(
        clk) );
  DFQD4BWP cu1_controlBlock_config__udcInit_0_reg_1_ ( .D(n332), .CP(
        cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu0_controlBlock_config__udcInit_0_reg_1_ ( .D(reset), .CP(
        cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu1_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(reset), 
        .CP(cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu1_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(n332), 
        .CP(cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu0_controlBlock_decXbar_config__outSelect_1_reg_0_ ( .D(n332), 
        .CP(cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu0_controlBlock_incXbar_config__outSelect_3_reg_1_ ( .D(n332), 
        .CP(cu0_controlBlock_incXbar_net4499) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_1_net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_1_net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_1_net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_1_net4403), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_1_net4400), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_1_net4397), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_FF_1_ff_reg_6_ ( .D(n123), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4412), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4409), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4406), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4403), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4400), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4397), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4394), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_4_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_4_net4391), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4412), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4409), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4406), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4403), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4400), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4397), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4394), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_5_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_5_net4391), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_1_net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_1_net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_2_ ( .D(
        cu1_RegisterBlock_FF_1_net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_1_net4403), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_1_net4400), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_1_net4397), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_6_ ( .D(
        cu1_RegisterBlock_FF_1_net4394), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_FF_1_ff_reg_7_ ( .D(n122), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4412), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4409), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4406), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4403), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4400), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4397), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_5_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_5_net4394), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4412), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4409), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4406), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4403), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4400), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4397), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4394), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_4_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_4_net4391), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_2_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_2_net4412), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_2_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_2_net4409), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_2_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_2_net4406), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4412), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4409), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4406), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4403), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4400), .CP(clk) );
  DFQD4BWP cu0_RegisterBlock_1_FF_3_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_3_net4397), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_2_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_2_net4412), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_2_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_2_net4409), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_2_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_2_net4406), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4412), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4409), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4406), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4403), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4400), .CP(clk) );
  DFQD4BWP cu1_RegisterBlock_1_FF_3_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_3_net4397), .CP(clk) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_5_ ( .D(cu1_RegisterBlock_FF_1_net4397), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .D(
        cu0_counterChain_CounterRC_counter_reg__net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_0_out_2_) );
  DFQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_2_ ( .D(
        cu1_counterChain_CounterRC_counter_reg__net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_0_out_2_) );
  DFQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .D(
        cu1_counterChain_CounterRC_1_counter_reg__net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_1_out_0_) );
  DFQD1BWP controlBox_commandReg_reg ( .D(controlBox_N6), .CP(clk), .Q(
        controlBox_commandReg) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_4_net4412), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[0]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_4_net4409), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[1]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_4_net4406), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[2]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_4_net4403), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[3]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_4_net4400), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[4]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_4_net4397), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[5]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_6_ ( .D(
        cu0_RegisterBlock_FF_4_net4394), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[6]) );
  DFQD1BWP cu0_RegisterBlock_FF_4_ff_reg_7_ ( .D(
        cu0_RegisterBlock_FF_4_net4391), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_2[7]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_5_net4412), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[0]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_5_net4409), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[1]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_5_net4406), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[2]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_5_net4403), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[3]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_5_net4400), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[4]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_5_net4397), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[5]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_6_ ( .D(
        cu0_RegisterBlock_FF_5_net4394), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[6]) );
  DFQD1BWP cu0_RegisterBlock_FF_5_ff_reg_7_ ( .D(
        cu0_RegisterBlock_FF_5_net4391), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_3[7]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_4_net4412), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_4_net4409), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[1]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_2_ ( .D(
        cu1_RegisterBlock_FF_4_net4406), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[2]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_4_net4403), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[3]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_4_net4400), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[4]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_4_net4397), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[5]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_6_ ( .D(
        cu1_RegisterBlock_FF_4_net4394), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[6]) );
  DFQD1BWP cu1_RegisterBlock_FF_4_ff_reg_7_ ( .D(
        cu1_RegisterBlock_FF_4_net4391), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_2[7]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_5_net4412), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_5_net4409), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[1]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_2_ ( .D(
        cu1_RegisterBlock_FF_5_net4406), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[2]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_5_net4403), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[3]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_5_net4400), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[4]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_5_net4397), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[5]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_6_ ( .D(
        cu1_RegisterBlock_FF_5_net4394), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[6]) );
  DFQD1BWP cu1_RegisterBlock_FF_5_ff_reg_7_ ( .D(
        cu1_RegisterBlock_FF_5_net4391), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_3[7]) );
  DFQD1BWP cu0_RegisterBlock_FF_2_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_2_net4412), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[0]) );
  DFQD1BWP cu0_RegisterBlock_FF_2_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_2_net4409), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[1]) );
  DFQD1BWP cu0_RegisterBlock_FF_2_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_2_net4406), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_0[2]) );
  DFQD1BWP cu1_RegisterBlock_FF_2_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_2_net4412), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_2_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_2_net4409), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[1]) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4412), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_6_ ( .D(cu1_RegisterBlock_FF_1_net4394), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4412), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4409), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4406), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4403), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4400), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4397), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4394), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4409), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4406), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4403), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_3_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4400), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_4_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4397), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4394), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4391), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu1_RegisterBlock_1_FF_1_io_data_out_7_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_0_ ( .D(cu0_RegisterBlock_FF_1_net4412), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_1_ ( .D(cu0_RegisterBlock_FF_1_net4409), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_3_ ( .D(cu0_RegisterBlock_FF_1_net4403), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_6_ ( .D(n123), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_6_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_2_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_2_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_3_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4403), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_4_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4400), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_5_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4397), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_6_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4394), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_2_ ( .D(cu1_RegisterBlock_FF_1_net4406), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_4_ ( .D(cu1_RegisterBlock_FF_1_net4400), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_4_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_0_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_0_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_1_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_2_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_3_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4403), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_3_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_4_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4400), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_4_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_5_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4397), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_5_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_6_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4394), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_1_FF_io_data_out_6_) );
  DFQD1BWP cu1_RegisterBlock_1_FF_ff_reg_7_ ( .D(
        cu1_RegisterBlock_1_FF_1_net4391), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_1_ ( .D(
        cu0_RegisterBlock_FF_3_net4409), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[1]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_2_ ( .D(
        cu0_RegisterBlock_FF_3_net4406), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[2]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_3_ ( .D(
        cu0_RegisterBlock_FF_3_net4403), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[3]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_4_ ( .D(
        cu0_RegisterBlock_FF_3_net4400), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[4]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_5_ ( .D(
        cu0_RegisterBlock_FF_3_net4397), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[5]) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .D(
        cu1_controlBlock_UpDownCtr_1_reg__net4469), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .D(
        cu0_controlBlock_UpDownCtr_reg__net4469), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_3_ ( .D(
        cu0_controlBlock_UpDownCtr_1_reg__net4469), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_3_ ( .D(
        cu1_controlBlock_UpDownCtr_reg__net4469), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .D(
        cu1_controlBlock_UpDownCtr_1_reg__net4472), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .D(
        cu0_controlBlock_UpDownCtr_reg__net4472), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_2_ ( .D(
        cu0_controlBlock_UpDownCtr_1_reg__net4472), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_2_ ( .D(
        cu1_controlBlock_UpDownCtr_reg__net4472), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_3_ ( .D(cu1_RegisterBlock_FF_1_net4403), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_3_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_5_ ( .D(cu0_RegisterBlock_FF_1_net4397), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_5_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_4_ ( .D(cu0_RegisterBlock_FF_1_net4400), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_4_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_0_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_0_) );
  DFQD1BWP cu0_RegisterBlock_1_FF_ff_reg_1_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_1_FF_io_data_out_1_) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_1_ ( .D(
        cu1_RegisterBlock_FF_3_net4409), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[1]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_2_ ( .D(
        cu1_RegisterBlock_FF_3_net4406), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[2]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_3_ ( .D(
        cu1_RegisterBlock_FF_3_net4403), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[3]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_4_ ( .D(
        cu1_RegisterBlock_FF_3_net4400), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[4]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_5_ ( .D(
        cu1_RegisterBlock_FF_3_net4397), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[5]) );
  DFQD1BWP cu0_RegisterBlock_FF_3_ff_reg_0_ ( .D(
        cu0_RegisterBlock_FF_3_net4412), .CP(clk), .Q(
        cu0_RegisterBlock_io_passDataOut_1[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_3_ff_reg_0_ ( .D(
        cu1_RegisterBlock_FF_3_net4412), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_1[0]) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_1_ ( .D(cu1_RegisterBlock_FF_1_net4409), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_1_) );
  DFQD1BWP cu0_RegisterBlock_FF_ff_reg_2_ ( .D(cu0_RegisterBlock_FF_1_net4406), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_RegisterBlock_FF_io_data_out_2_) );
  DFQD1BWP cu1_RegisterBlock_FF_ff_reg_0_ ( .D(cu1_RegisterBlock_FF_1_net4412), 
        .CP(cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_RegisterBlock_FF_io_data_out_0_) );
  DFQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .D(
        cu0_counterChain_CounterRC_counter_reg__net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_0_out_1_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .D(
        cu1_controlBlock_UpDownCtr_1_reg__net4478), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .D(
        cu0_controlBlock_UpDownCtr_reg__net4478), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_0_ ( .D(
        cu0_controlBlock_UpDownCtr_1_reg__net4478), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_0_ ( .D(
        cu1_controlBlock_UpDownCtr_reg__net4478), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .D(
        cu1_controlBlock_UpDownCtr_1_reg__net4475), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .D(
        cu0_controlBlock_UpDownCtr_reg__net4475), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFQD1BWP cu0_controlBlock_UpDownCtr_1_reg__ff_reg_1_ ( .D(
        cu0_controlBlock_UpDownCtr_1_reg__net4475), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_) );
  DFQD1BWP cu1_controlBlock_UpDownCtr_reg__ff_reg_1_ ( .D(
        cu1_controlBlock_UpDownCtr_reg__net4475), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_) );
  DFQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .D(
        cu0_counterChain_CounterRC_1_counter_reg__net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_1_out_2_) );
  DFQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_2_ ( .D(
        cu1_counterChain_CounterRC_1_counter_reg__net4406), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_1_out_2_) );
  DFQD1BWP cu1_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .D(
        cu1_counterChain_CounterRC_1_counter_reg__net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_1_out_1_) );
  DFQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_1_ ( .D(
        cu0_counterChain_CounterRC_1_counter_reg__net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_1_out_1_) );
  DFQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_1_ ( .D(
        cu1_counterChain_CounterRC_counter_reg__net4409), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_0_out_1_) );
  DFQD1BWP cu0_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .D(
        cu0_counterChain_CounterRC_counter_reg__net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_0_out_0_) );
  DFQD1BWP cu1_counterChain_CounterRC_counter_reg__ff_reg_0_ ( .D(
        cu1_counterChain_CounterRC_counter_reg__net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_io_data_0_out_0_) );
  DFQD1BWP cu0_counterChain_CounterRC_1_counter_reg__ff_reg_0_ ( .D(
        cu0_counterChain_CounterRC_1_counter_reg__net4412), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu0_counterChain_io_data_1_out_0_) );
  DFQD1BWP cu1_counterChain_CounterRC_config__stride_reg_0_ ( .D(n332), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415), .Q(
        cu1_counterChain_CounterRC_config__stride_0_) );
  DFQD2BWP cu1_RegisterBlock_FF_ff_reg_7_ ( .D(n122), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD2BWP cu0_RegisterBlock_FF_ff_reg_7_ ( .D(n118), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD2BWP cu0_RegisterBlock_1_FF_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4391), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFQD2BWP cu0_RegisterBlock_FF_1_ff_reg_7_ ( .D(n118), .CP(
        cu1_counterChain_CounterRC_1_counter_reg__net4415) );
  DFKCNQD1BWP cu1_RegisterBlock_1_FF_5_ff_reg_7_ ( .CN(n333), .D(
        cu1_RegisterBlock_io_passDataOut_3[7]), .CP(clk) );
  DFKCNQD1BWP cu1_RegisterBlock_FF_2_ff_reg_2_ ( .CN(n333), .D(
        cu1_counterChain_io_data_0_out_2_), .CP(clk), .Q(
        cu1_RegisterBlock_io_passDataOut_0[2]) );
  DFQD1BWP cu0_RegisterBlock_1_FF_1_ff_reg_7_ ( .D(
        cu0_RegisterBlock_1_FF_1_net4391), .CP(
        cu1_RegisterBlock_1_FF_1_net4415), .Q(
        cu0_RegisterBlock_1_FF_1_io_data_out_7_) );
  XNR2D1BWP U384 ( .A1(n271), .A2(n270), .ZN(cu1_IntFU_1_m_T3[7]) );
  INVD1BWP U385 ( .I(n236), .ZN(n197) );
  INVD1BWP U386 ( .I(n237), .ZN(n201) );
  IND2D1BWP U387 ( .A1(n191), .B1(n290), .ZN(n200) );
  INVD1BWP U388 ( .I(cu1_RegisterBlock_FF_io_data_out_0_), .ZN(n191) );
  INVD1BWP U389 ( .I(n229), .ZN(n202) );
  INVD1BWP U390 ( .I(n230), .ZN(n203) );
  INVD1BWP U391 ( .I(n244), .ZN(n176) );
  INVD1BWP U392 ( .I(n245), .ZN(n173) );
  ND2D1BWP U393 ( .A1(n290), .A2(cu0_RegisterBlock_FF_io_data_out_0_), .ZN(
        n157) );
  ND2D1BWP U394 ( .A1(n290), .A2(cu0_RegisterBlock_FF_io_data_out_1_), .ZN(
        n172) );
  INVD1BWP U395 ( .I(n256), .ZN(n179) );
  INVD1BWP U396 ( .I(n255), .ZN(n178) );
  ND2D1BWP U397 ( .A1(n290), .A2(cu0_RegisterBlock_FF_io_data_out_2_), .ZN(
        n171) );
  INVD1BWP U398 ( .I(n214), .ZN(n180) );
  INVD1BWP U399 ( .I(n215), .ZN(n177) );
  IOA21D1BWP U400 ( .A1(n294), .A2(cu0_counterChain_io_data_0_out_2_), .B(n171), .ZN(n244) );
  IOA21D1BWP U401 ( .A1(cu0_counterChain_io_data_1_out_2_), .A2(n268), .B(n171), .ZN(n245) );
  ND2D1BWP U402 ( .A1(n294), .A2(cu1_counterChain_io_data_0_out_0_), .ZN(n192)
         );
  IOA21D1BWP U403 ( .A1(cu1_counterChain_io_data_1_out_1_), .A2(n268), .B(n190), .ZN(n230) );
  ND2D1BWP U404 ( .A1(n196), .A2(n195), .ZN(n229) );
  ND2D1BWP U405 ( .A1(n194), .A2(n193), .ZN(n236) );
  ND2D1BWP U406 ( .A1(n194), .A2(n189), .ZN(n237) );
  INR2D1BWP U407 ( .A1(n294), .B1(n332), .ZN(n285) );
  INR2D1BWP U408 ( .A1(n333), .B1(n294), .ZN(n298) );
  FICOND1BWP U409 ( .A(n164), .B(n163), .CI(n162), .CON(n253), .S(
        cu0_IntFU_1_m_T3[4]) );
  IOA21D1BWP U410 ( .A1(n294), .A2(cu0_counterChain_io_data_1_out_1_), .B(n172), .ZN(n256) );
  CKND1BWP U411 ( .I(n233), .ZN(n93) );
  CKND1BWP U412 ( .I(n238), .ZN(n94) );
  AOI31D1BWP U413 ( .A1(n232), .A2(n239), .A3(n93), .B(n94), .ZN(n222) );
  AN3D1BWP U414 ( .A1(n290), .A2(n298), .A3(
        cu0_RegisterBlock_FF_io_data_out_6_), .Z(n118) );
  INR2D1BWP U415 ( .A1(n286), .B1(n289), .ZN(cu0_RegisterBlock_FF_3_net4403)
         );
  INR2D1BWP U416 ( .A1(cu1_IntFU_1_m_T3[5]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4397) );
  XNR3D1BWP U417 ( .A1(n253), .A2(n252), .A3(n251), .ZN(cu0_IntFU_1_m_T3[5])
         );
  CKND1BWP U418 ( .I(cu0_counterChain_io_data_0_out_1_), .ZN(n95) );
  OAI21D1BWP U419 ( .A1(n290), .A2(n95), .B(n172), .ZN(n255) );
  CKND1BWP U420 ( .I(n200), .ZN(n96) );
  AOI21D1BWP U421 ( .A1(n294), .A2(cu1_counterChain_io_data_1_out_0_), .B(n96), 
        .ZN(n119) );
  IND2D1BWP U422 ( .A1(n220), .B1(n221), .ZN(n97) );
  CKXOR2D1BWP U423 ( .A1(n222), .A2(n97), .Z(n288) );
  INR2D1BWP U424 ( .A1(cu1_IntFU_1_m_T3[6]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4394) );
  INR2D1BWP U425 ( .A1(cu1_IntFU_1_m_T3[4]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4400) );
  INR2D1BWP U426 ( .A1(cu1_IntFU_1_m_T3[3]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4403) );
  INR2D1BWP U427 ( .A1(cu0_IntFU_1_m_T3[5]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4397) );
  CKND1BWP U428 ( .I(n297), .ZN(n98) );
  AO31D1BWP U429 ( .A1(n290), .A2(n298), .A3(
        cu1_RegisterBlock_FF_io_data_out_4_), .B(n98), .Z(
        cu1_RegisterBlock_FF_1_net4397) );
  CKND2D1BWP U430 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_7_), .A2(n268), 
        .ZN(n99) );
  CKXOR2D1BWP U431 ( .A1(n99), .A2(n136), .Z(cu0_IntFU_1_m_T3[7]) );
  AN2D1BWP U432 ( .A1(n187), .A2(n186), .Z(n188) );
  INR2D1BWP U433 ( .A1(n232), .B1(n233), .ZN(n240) );
  IND3D1BWP U434 ( .A1(cu0_counterChain_io_data_1_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n333), .ZN(n326) );
  ND2D1BWP U435 ( .A1(n215), .A2(n214), .ZN(n254) );
  IND2D1BWP U436 ( .A1(n216), .B1(n217), .ZN(n100) );
  CKXOR2D1BWP U437 ( .A1(n218), .A2(n100), .Z(n286) );
  INR2D1BWP U438 ( .A1(cu0_IntFU_1_m_T3[6]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4394) );
  INR2D1BWP U439 ( .A1(cu0_IntFU_1_m_T3[4]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4400) );
  INR2D1BWP U440 ( .A1(cu0_IntFU_1_m_T3[1]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4409) );
  CKND2D1BWP U441 ( .A1(cu1_RegisterBlock_FF_io_data_out_3_), .A2(n298), .ZN(
        n101) );
  OAI21D1BWP U442 ( .A1(n101), .A2(n294), .B(n295), .ZN(
        cu1_RegisterBlock_FF_1_net4400) );
  AN2D1BWP U443 ( .A1(n151), .A2(n152), .Z(n102) );
  CKND1BWP U444 ( .I(n152), .ZN(n103) );
  AOI21D1BWP U445 ( .A1(cu1_RegisterBlock_1_FF_1_io_data_out_3_), .A2(n294), 
        .B(n103), .ZN(n104) );
  MAOI222D1BWP U446 ( .A(n170), .B(n102), .C(n104), .ZN(n159) );
  XNR3D1BWP U447 ( .A1(n170), .A2(n102), .A3(n104), .ZN(cu1_IntFU_1_m_T3[3])
         );
  CKND2D1BWP U448 ( .A1(n290), .A2(cu1_RegisterBlock_FF_io_data_out_2_), .ZN(
        n194) );
  IND3D1BWP U449 ( .A1(cu1_counterChain_io_data_0_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n333), .ZN(n328) );
  OA21D1BWP U450 ( .A1(n258), .A2(n257), .B(n259), .Z(n281) );
  CKND1BWP U451 ( .I(n291), .ZN(n219) );
  AN2D1BWP U452 ( .A1(n290), .A2(cu0_RegisterBlock_FF_io_data_out_3_), .Z(n293) );
  IAO21D1BWP U453 ( .A1(n231), .A2(n232), .B(n240), .ZN(n282) );
  INR2D1BWP U454 ( .A1(cu0_IntFU_1_m_T3[7]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4391) );
  INR2D1BWP U455 ( .A1(n288), .B1(n289), .ZN(cu1_RegisterBlock_FF_3_net4403)
         );
  INR2D1BWP U456 ( .A1(cu1_IntFU_1_m_T3[2]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4406) );
  INR2D1BWP U457 ( .A1(cu1_IntFU_1_m_T3[1]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4409) );
  INR2D1BWP U458 ( .A1(cu1_IntFU_1_m_T3[0]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_1_net4412) );
  INR2D1BWP U459 ( .A1(cu1_RegisterBlock_io_passDataOut_1[0]), .B1(n332), .ZN(
        cu1_RegisterBlock_1_FF_3_net4412) );
  AN3D1BWP U460 ( .A1(n290), .A2(n298), .A3(
        cu0_RegisterBlock_FF_io_data_out_5_), .Z(n123) );
  OA21D1BWP U461 ( .A1(n290), .A2(n301), .B(n129), .Z(n105) );
  CKND1BWP U462 ( .I(n129), .ZN(n106) );
  AOI21D1BWP U463 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_3_), .A2(n294), 
        .B(n106), .ZN(n107) );
  MAOI222D1BWP U464 ( .A(n169), .B(n105), .C(n107), .ZN(n162) );
  XNR3D1BWP U465 ( .A1(n169), .A2(n105), .A3(n107), .ZN(cu0_IntFU_1_m_T3[3])
         );
  AN2D1BWP U466 ( .A1(n147), .A2(n148), .Z(n108) );
  CKND1BWP U467 ( .I(n148), .ZN(n109) );
  AOI21D1BWP U468 ( .A1(n268), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_5_), 
        .B(n109), .ZN(n110) );
  MAOI222D1BWP U469 ( .A(n168), .B(n108), .C(n110), .ZN(n269) );
  XNR3D1BWP U470 ( .A1(n168), .A2(n108), .A3(n110), .ZN(cu1_IntFU_1_m_T3[5])
         );
  AN2D1BWP U471 ( .A1(n206), .A2(n207), .Z(n121) );
  IND3D1BWP U472 ( .A1(cu1_counterChain_io_data_1_out_2_), .B1(
        cu1_counterChain_CounterRC_config__stride_0_), .B2(n333), .ZN(n330) );
  INR2D1BWP U473 ( .A1(cu0_IntFU_1_m_T3[3]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4403) );
  INR2D1BWP U474 ( .A1(cu0_IntFU_1_m_T3[2]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4406) );
  INR2D1BWP U475 ( .A1(cu0_IntFU_1_m_T3[0]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_1_net4412) );
  INR2D1BWP U476 ( .A1(cu1_counterChain_io_data_0_out_1_), .B1(n332), .ZN(
        cu1_RegisterBlock_FF_2_net4409) );
  INR2D1BWP U477 ( .A1(cu1_counterChain_io_data_0_out_0_), .B1(n332), .ZN(
        cu1_RegisterBlock_FF_2_net4412) );
  INR2D1BWP U478 ( .A1(cu0_counterChain_io_data_0_out_1_), .B1(n332), .ZN(
        cu0_RegisterBlock_FF_2_net4409) );
  INR2D1BWP U479 ( .A1(cu0_counterChain_io_data_0_out_0_), .B1(n332), .ZN(
        cu0_RegisterBlock_FF_2_net4412) );
  INR2D1BWP U480 ( .A1(cu1_RegisterBlock_io_passDataOut_1[5]), .B1(reset), 
        .ZN(cu1_RegisterBlock_1_FF_3_net4397) );
  INR2D1BWP U481 ( .A1(cu1_RegisterBlock_io_passDataOut_1[4]), .B1(reset), 
        .ZN(cu1_RegisterBlock_1_FF_3_net4400) );
  INR2D1BWP U482 ( .A1(cu1_RegisterBlock_io_passDataOut_1[3]), .B1(reset), 
        .ZN(cu1_RegisterBlock_1_FF_3_net4403) );
  INR2D1BWP U483 ( .A1(cu1_RegisterBlock_io_passDataOut_1[2]), .B1(reset), 
        .ZN(cu1_RegisterBlock_1_FF_3_net4406) );
  INR2D1BWP U484 ( .A1(cu1_RegisterBlock_io_passDataOut_1[1]), .B1(reset), 
        .ZN(cu1_RegisterBlock_1_FF_3_net4409) );
  INR2D1BWP U485 ( .A1(cu0_RegisterBlock_io_passDataOut_1[0]), .B1(n332), .ZN(
        cu0_RegisterBlock_1_FF_3_net4412) );
  INR2D1BWP U486 ( .A1(cu1_mem0raMux_io_out_0[3]), .B1(reset), .ZN(
        cu1_RegisterBlock_FF_1_net4403) );
  INR2D1BWP U487 ( .A1(cu1_mem0raMux_io_out_0[1]), .B1(n332), .ZN(
        cu1_RegisterBlock_FF_1_net4409) );
  INR2D1BWP U488 ( .A1(cu1_mem0raMux_io_out_0[0]), .B1(n332), .ZN(
        cu1_RegisterBlock_FF_1_net4412) );
  CKND1BWP U489 ( .I(n296), .ZN(n111) );
  AO31D1BWP U490 ( .A1(n290), .A2(n298), .A3(
        cu0_RegisterBlock_FF_io_data_out_4_), .B(n111), .Z(
        cu0_RegisterBlock_FF_1_net4397) );
  INR2D1BWP U491 ( .A1(cu0_mem1raMux_io_out_0[3]), .B1(n332), .ZN(
        cu0_RegisterBlock_FF_1_net4403) );
  INR2D1BWP U492 ( .A1(cu0_mem1raMux_io_out_0[2]), .B1(reset), .ZN(
        cu0_RegisterBlock_FF_1_net4406) );
  INR2D1BWP U493 ( .A1(cu0_mem1raMux_io_out_0[1]), .B1(n332), .ZN(
        cu0_RegisterBlock_FF_1_net4409) );
  CKND1BWP U494 ( .I(n127), .ZN(n112) );
  AOI31D1BWP U495 ( .A1(n156), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_6_), 
        .A3(n294), .B(n112), .ZN(n136) );
  ND3D1BWP U496 ( .A1(cu0_RegisterBlock_1_FF_1_io_data_out_6_), .A2(n294), 
        .A3(n127), .ZN(n113) );
  XNR2D1BWP U497 ( .A1(n113), .A2(n156), .ZN(cu0_IntFU_1_m_T3[6]) );
  IOA21D1BWP U498 ( .A1(n268), .A2(cu1_RegisterBlock_io_passDataOut_1[0]), .B(
        n139), .ZN(n114) );
  IOA21D1BWP U499 ( .A1(n294), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_0_), 
        .B(n139), .ZN(n115) );
  CKND2D1BWP U500 ( .A1(n114), .A2(n115), .ZN(n165) );
  CKXOR2D1BWP U501 ( .A1(n114), .A2(n115), .Z(cu1_IntFU_1_m_T3[0]) );
  CKND1BWP U502 ( .I(n146), .ZN(n116) );
  AOI31D1BWP U503 ( .A1(n269), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_6_), 
        .A3(n294), .B(n116), .ZN(n270) );
  ND3D1BWP U504 ( .A1(cu1_RegisterBlock_1_FF_1_io_data_out_6_), .A2(n294), 
        .A3(n146), .ZN(n117) );
  XNR2D1BWP U505 ( .A1(n117), .A2(n269), .ZN(cu1_IntFU_1_m_T3[6]) );
  BUFFD4BWP U506 ( .I(cu0_T21_0_), .Z(n294) );
  INVD6BWP U507 ( .I(cu0_T21_0_), .ZN(n290) );
  AO21D1BWP U508 ( .A1(n226), .A2(n225), .B(n188), .Z(n120) );
  AN2XD1BWP U509 ( .A1(n267), .A2(n298), .Z(n122) );
  AO21D1BWP U510 ( .A1(n213), .A2(n212), .B(n121), .Z(n124) );
  BUFFD2BWP U511 ( .I(cu0_T21_0_), .Z(n268) );
  AN2XD1BWP U512 ( .A1(n200), .A2(n192), .Z(n125) );
  CKND2BWP U513 ( .I(reset), .ZN(n333) );
  INVD1BWP U514 ( .I(n333), .ZN(n332) );
  XOR2D1BWP U515 ( .A1(n206), .A2(n207), .Z(n209) );
  XOR2D1BWP U516 ( .A1(n186), .A2(n187), .Z(n185) );
  INR2D1BWP U517 ( .A1(cu1_RegisterBlock_FF_io_data_out_5_), .B1(n268), .ZN(
        n126) );
  AN2D1BWP U518 ( .A1(n298), .A2(n126), .Z(cu1_RegisterBlock_FF_1_net4394) );
  ND2D1BWP U519 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_6_), .ZN(
        n127) );
  ND2D1BWP U520 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_4_), .ZN(
        n128) );
  IOA21D1BWP U521 ( .A1(n294), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_4_), 
        .B(n128), .ZN(n164) );
  CKND1BWP U522 ( .I(cu0_RegisterBlock_io_passDataOut_1[4]), .ZN(n302) );
  OAI21D1BWP U523 ( .A1(n290), .A2(n302), .B(n128), .ZN(n163) );
  ND2D1BWP U524 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_3_), .ZN(
        n129) );
  CKND1BWP U525 ( .I(cu0_RegisterBlock_io_passDataOut_1[3]), .ZN(n301) );
  ND2D1BWP U526 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_1_), .ZN(
        n130) );
  IOA21D1BWP U527 ( .A1(n268), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_1_), 
        .B(n130), .ZN(n145) );
  CKND1BWP U528 ( .I(cu0_RegisterBlock_io_passDataOut_1[1]), .ZN(n299) );
  OAI21D1BWP U529 ( .A1(n290), .A2(n299), .B(n130), .ZN(n144) );
  ND2D1BWP U530 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_0_), .ZN(
        n131) );
  IOA21D1BWP U531 ( .A1(n294), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_0_), 
        .B(n131), .ZN(n266) );
  IOA21D1BWP U532 ( .A1(n268), .A2(cu0_RegisterBlock_io_passDataOut_1[0]), .B(
        n131), .ZN(n265) );
  CKND1BWP U533 ( .I(cu0_RegisterBlock_io_passDataOut_1[2]), .ZN(n300) );
  ND2D1BWP U534 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_2_), .ZN(
        n132) );
  OAI21D1BWP U535 ( .A1(n290), .A2(n300), .B(n132), .ZN(n262) );
  IOA21D1BWP U536 ( .A1(n268), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_2_), 
        .B(n132), .ZN(n261) );
  AN2XD1BWP U537 ( .A1(n262), .A2(n261), .Z(n133) );
  OAI22D1BWP U538 ( .A1(n264), .A2(n133), .B1(n262), .B2(n261), .ZN(n169) );
  CKND1BWP U539 ( .I(cu0_RegisterBlock_io_passDataOut_1[5]), .ZN(n303) );
  ND2D1BWP U540 ( .A1(n290), .A2(cu0_RegisterBlock_1_FF_io_data_out_5_), .ZN(
        n134) );
  OAI21D1BWP U541 ( .A1(n290), .A2(n303), .B(n134), .ZN(n252) );
  IOA21D1BWP U542 ( .A1(n268), .A2(cu0_RegisterBlock_1_FF_1_io_data_out_5_), 
        .B(n134), .ZN(n251) );
  NR2D1BWP U543 ( .A1(n252), .A2(n251), .ZN(n135) );
  MOAI22D1BWP U544 ( .A1(n253), .A2(n135), .B1(n251), .B2(n252), .ZN(n156) );
  ND2D1BWP U545 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_2_), .ZN(
        n138) );
  IOA21D1BWP U546 ( .A1(n294), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_2_), 
        .B(n138), .ZN(n155) );
  CKND2D1BWP U547 ( .A1(n268), .A2(cu1_RegisterBlock_io_passDataOut_1[2]), 
        .ZN(n137) );
  ND2D1BWP U548 ( .A1(n138), .A2(n137), .ZN(n154) );
  ND2D1BWP U549 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_0_), .ZN(
        n139) );
  ND2D1BWP U550 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_1_), .ZN(
        n141) );
  CKND2D1BWP U551 ( .A1(n268), .A2(cu1_RegisterBlock_io_passDataOut_1[1]), 
        .ZN(n140) );
  ND2D1BWP U552 ( .A1(n141), .A2(n140), .ZN(n166) );
  IOA21D1BWP U553 ( .A1(n294), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_1_), 
        .B(n141), .ZN(n167) );
  NR2D1BWP U554 ( .A1(n166), .A2(n167), .ZN(n142) );
  MOAI22D1BWP U555 ( .A1(n165), .A2(n142), .B1(n167), .B2(n166), .ZN(n153) );
  FICIND2BWP U556 ( .CIN(n143), .B(n144), .A(n145), .CO(n264), .S(
        cu0_IntFU_1_m_T3[1]) );
  ND2D1BWP U557 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_6_), .ZN(
        n146) );
  ND2D1BWP U558 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_5_), .ZN(
        n148) );
  CKND2D1BWP U559 ( .A1(n294), .A2(cu1_RegisterBlock_io_passDataOut_1[5]), 
        .ZN(n147) );
  ND2D1BWP U560 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_4_), .ZN(
        n150) );
  IOA21D1BWP U561 ( .A1(n294), .A2(cu1_RegisterBlock_1_FF_1_io_data_out_4_), 
        .B(n150), .ZN(n161) );
  CKND2D1BWP U562 ( .A1(n268), .A2(cu1_RegisterBlock_io_passDataOut_1[4]), 
        .ZN(n149) );
  ND2D1BWP U563 ( .A1(n150), .A2(n149), .ZN(n160) );
  ND2D1BWP U564 ( .A1(n290), .A2(cu1_RegisterBlock_1_FF_io_data_out_3_), .ZN(
        n152) );
  CKND2D1BWP U565 ( .A1(n268), .A2(cu1_RegisterBlock_io_passDataOut_1[3]), 
        .ZN(n151) );
  FICOND1BWP U566 ( .A(n155), .B(n154), .CI(n153), .CON(n170), .S(
        cu1_IntFU_1_m_T3[2]) );
  IOA21D1BWP U567 ( .A1(n294), .A2(cu0_counterChain_io_data_0_out_0_), .B(n157), .ZN(n214) );
  CKND1BWP U568 ( .I(cu0_counterChain_io_data_1_out_0_), .ZN(n158) );
  OAI21D1BWP U569 ( .A1(n158), .A2(n290), .B(n157), .ZN(n215) );
  NR2D1BWP U570 ( .A1(n180), .A2(n177), .ZN(n278) );
  AN2D1BWP U571 ( .A1(n268), .A2(n278), .Z(cu0_mem1raMux_io_out_0[0]) );
  FICOND2BWP U572 ( .A(n161), .B(n160), .CI(n159), .CON(n168), .S(
        cu1_IntFU_1_m_T3[4]) );
  XNR3D1BWP U573 ( .A1(n167), .A2(n166), .A3(n165), .ZN(cu1_IntFU_1_m_T3[1])
         );
  NR2D1BWP U574 ( .A1(n176), .A2(n179), .ZN(n187) );
  NR2D1BWP U575 ( .A1(n180), .A2(n173), .ZN(n175) );
  NR2D1BWP U576 ( .A1(n178), .A2(n179), .ZN(n174) );
  NR2D1BWP U577 ( .A1(n178), .A2(n173), .ZN(n184) );
  NR2D1BWP U578 ( .A1(n185), .A2(n184), .ZN(n216) );
  HA1D1BWP U579 ( .A(n175), .B(n174), .CO(n186), .S(n182) );
  NR2D1BWP U580 ( .A1(n176), .A2(n177), .ZN(n181) );
  OR2XD1BWP U581 ( .A1(n182), .A2(n181), .Z(n247) );
  NR2D1BWP U582 ( .A1(n178), .A2(n177), .ZN(n258) );
  NR2D1BWP U583 ( .A1(n180), .A2(n179), .ZN(n257) );
  ND2D1BWP U584 ( .A1(n258), .A2(n257), .ZN(n259) );
  CKND1BWP U585 ( .I(n259), .ZN(n248) );
  ND2D1BWP U586 ( .A1(n182), .A2(n181), .ZN(n246) );
  CKND1BWP U587 ( .I(n246), .ZN(n183) );
  AOI21D1BWP U588 ( .A1(n247), .A2(n248), .B(n183), .ZN(n218) );
  ND2D1BWP U589 ( .A1(n185), .A2(n184), .ZN(n217) );
  OAI21D1BWP U590 ( .A1(n216), .A2(n218), .B(n217), .ZN(n226) );
  AN2XD1BWP U591 ( .A1(n244), .A2(n245), .Z(n225) );
  CKND1BWP U592 ( .I(n188), .ZN(n224) );
  ND2D1BWP U593 ( .A1(n120), .A2(n285), .ZN(n296) );
  CKND1BWP U594 ( .I(n296), .ZN(cu0_RegisterBlock_FF_3_net4397) );
  ND2D1BWP U595 ( .A1(n268), .A2(cu1_counterChain_io_data_0_out_2_), .ZN(n189)
         );
  IND2D1BWP U596 ( .A1(cu0_T21_0_), .B1(cu1_RegisterBlock_FF_io_data_out_1_), 
        .ZN(n190) );
  NR2D1BWP U597 ( .A1(n201), .A2(n203), .ZN(n207) );
  ND2D1BWP U598 ( .A1(n268), .A2(cu1_counterChain_io_data_1_out_2_), .ZN(n193)
         );
  NR2D1BWP U599 ( .A1(n125), .A2(n197), .ZN(n199) );
  ND2D1BWP U600 ( .A1(n290), .A2(cu1_RegisterBlock_FF_io_data_out_1_), .ZN(
        n196) );
  ND2D1BWP U601 ( .A1(n294), .A2(cu1_counterChain_io_data_0_out_1_), .ZN(n195)
         );
  NR2D1BWP U602 ( .A1(n202), .A2(n203), .ZN(n198) );
  NR2D1BWP U603 ( .A1(n202), .A2(n197), .ZN(n208) );
  NR2D1BWP U604 ( .A1(n201), .A2(n197), .ZN(n212) );
  IND2D1BWP U605 ( .A1(n121), .B1(n212), .ZN(n210) );
  HA1D1BWP U606 ( .A(n199), .B(n198), .CO(n206), .S(n205) );
  NR2D1BWP U607 ( .A1(n201), .A2(n119), .ZN(n204) );
  OR2XD1BWP U608 ( .A1(n205), .A2(n204), .Z(n239) );
  NR2D1BWP U609 ( .A1(n202), .A2(n119), .ZN(n231) );
  CKND1BWP U610 ( .I(n231), .ZN(n233) );
  NR2D1BWP U611 ( .A1(n125), .A2(n203), .ZN(n232) );
  ND2D1BWP U612 ( .A1(n205), .A2(n204), .ZN(n238) );
  NR2D1BWP U613 ( .A1(n209), .A2(n208), .ZN(n220) );
  ND2D1BWP U614 ( .A1(n209), .A2(n208), .ZN(n221) );
  OAI21D1BWP U615 ( .A1(n222), .A2(n220), .B(n221), .ZN(n213) );
  XNR2D1BWP U616 ( .A1(n210), .A2(n213), .ZN(n211) );
  ND2D1BWP U617 ( .A1(n211), .A2(n285), .ZN(n295) );
  CKND1BWP U618 ( .I(n295), .ZN(cu1_RegisterBlock_FF_3_net4400) );
  ND2D1BWP U619 ( .A1(n124), .A2(n285), .ZN(n297) );
  CKND1BWP U620 ( .I(n297), .ZN(cu1_RegisterBlock_FF_3_net4397) );
  MUX2D1BWP U621 ( .I0(n219), .I1(n286), .S(n294), .Z(
        cu0_mem1raMux_io_out_0[3]) );
  MUX2D1BWP U622 ( .I0(n223), .I1(n288), .S(n294), .Z(
        cu1_mem0raMux_io_out_0[3]) );
  ND2D1BWP U623 ( .A1(n225), .A2(n224), .ZN(n227) );
  XNR2D1BWP U624 ( .A1(n227), .A2(n226), .ZN(n228) );
  ND2D1BWP U625 ( .A1(n228), .A2(n285), .ZN(n292) );
  CKND1BWP U626 ( .I(n292), .ZN(cu0_RegisterBlock_FF_3_net4400) );
  FICIND1BWP U627 ( .CIN(n119), .B(n229), .A(n230), .CO(n235), .S(n234) );
  MUX2D1BWP U628 ( .I0(n234), .I1(n282), .S(n294), .Z(
        cu1_mem0raMux_io_out_0[1]) );
  FA1D1BWP U629 ( .A(n237), .B(n236), .CI(n235), .CO(n223), .S(n242) );
  ND2D1BWP U630 ( .A1(n239), .A2(n238), .ZN(n241) );
  XNR2D1BWP U631 ( .A1(n241), .A2(n240), .ZN(n283) );
  MUX2D1BWP U632 ( .I0(n242), .I1(n283), .S(n268), .Z(
        cu1_mem0raMux_io_out_0[2]) );
  FICOND1BWP U633 ( .A(n245), .B(n244), .CI(n243), .CON(n291), .S(n250) );
  ND2D1BWP U634 ( .A1(n247), .A2(n246), .ZN(n249) );
  XNR2D1BWP U635 ( .A1(n249), .A2(n248), .ZN(n284) );
  MUX2D1BWP U636 ( .I0(n250), .I1(n284), .S(n294), .Z(
        cu0_mem1raMux_io_out_0[2]) );
  NR2D1BWP U637 ( .A1(n125), .A2(n119), .ZN(n279) );
  AN2D1BWP U638 ( .A1(n294), .A2(n279), .Z(cu1_mem0raMux_io_out_0[0]) );
  FICIND1BWP U639 ( .CIN(n254), .B(n255), .A(n256), .CO(n243), .S(n260) );
  MUX2D1BWP U640 ( .I0(n260), .I1(n281), .S(n294), .Z(
        cu0_mem1raMux_io_out_0[1]) );
  XOR2D1BWP U641 ( .A1(n262), .A2(n261), .Z(n263) );
  XOR2D1BWP U642 ( .A1(n264), .A2(n263), .Z(cu0_IntFU_1_m_T3[2]) );
  HICOND1BWP U643 ( .A(n266), .CI(n265), .CON(n143), .S(cu0_IntFU_1_m_T3[0])
         );
  CKND1BWP U644 ( .I(n298), .ZN(cu1_RegisterBlock_1_FF_1_net4388) );
  AN2XD1BWP U645 ( .A1(controlBox_commandReg), .A2(n333), .Z(
        controlBox_pulser_N3) );
  AN2XD1BWP U646 ( .A1(cu1_RegisterBlock_io_passDataOut_2[4]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4400) );
  AN2XD1BWP U647 ( .A1(cu1_RegisterBlock_io_passDataOut_2[3]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4403) );
  AN2XD1BWP U648 ( .A1(cu1_RegisterBlock_io_passDataOut_2[2]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4406) );
  AN2XD1BWP U649 ( .A1(cu1_RegisterBlock_io_passDataOut_2[1]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4409) );
  AN2XD1BWP U650 ( .A1(cu0_RegisterBlock_io_passDataOut_2[4]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4400) );
  AN2XD1BWP U651 ( .A1(cu1_RegisterBlock_io_passDataOut_2[0]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4412) );
  AN2XD1BWP U652 ( .A1(cu0_RegisterBlock_io_passDataOut_2[7]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4391) );
  AN2XD1BWP U653 ( .A1(cu0_RegisterBlock_io_passDataOut_3[1]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4409) );
  AN2XD1BWP U654 ( .A1(cu0_RegisterBlock_io_passDataOut_3[5]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4397) );
  AN2XD1BWP U655 ( .A1(cu0_RegisterBlock_io_passDataOut_3[7]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4391) );
  AN2XD1BWP U656 ( .A1(cu0_RegisterBlock_io_passDataOut_2[0]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4412) );
  AN2XD1BWP U657 ( .A1(cu0_RegisterBlock_io_passDataOut_0[1]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_2_net4409) );
  AN2XD1BWP U658 ( .A1(cu1_RegisterBlock_io_passDataOut_2[7]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4391) );
  AN2XD1BWP U659 ( .A1(cu1_RegisterBlock_io_passDataOut_0[0]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_2_net4412) );
  AN2XD1BWP U660 ( .A1(cu1_RegisterBlock_io_passDataOut_0[2]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_2_net4406) );
  AN2XD1BWP U661 ( .A1(cu1_RegisterBlock_io_passDataOut_0[1]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_2_net4409) );
  AN2XD1BWP U662 ( .A1(cu1_RegisterBlock_io_passDataOut_2[6]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4394) );
  AN2XD1BWP U663 ( .A1(cu1_RegisterBlock_io_passDataOut_2[5]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_4_net4397) );
  AN2XD1BWP U664 ( .A1(cu1_RegisterBlock_io_passDataOut_3[0]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4412) );
  AN2XD1BWP U665 ( .A1(cu1_RegisterBlock_io_passDataOut_3[1]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4409) );
  AN2XD1BWP U666 ( .A1(cu1_RegisterBlock_io_passDataOut_3[2]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4406) );
  AN2XD1BWP U667 ( .A1(cu1_RegisterBlock_io_passDataOut_3[3]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4403) );
  AN2XD1BWP U668 ( .A1(cu0_RegisterBlock_io_passDataOut_0[2]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_2_net4406) );
  AN2XD1BWP U669 ( .A1(cu1_RegisterBlock_io_passDataOut_3[4]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4400) );
  AN2XD1BWP U670 ( .A1(cu1_RegisterBlock_io_passDataOut_3[5]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4397) );
  AN2XD1BWP U671 ( .A1(cu1_RegisterBlock_io_passDataOut_3[6]), .A2(n333), .Z(
        cu1_RegisterBlock_1_FF_5_net4394) );
  AN2XD1BWP U672 ( .A1(cu0_RegisterBlock_io_passDataOut_0[0]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_2_net4412) );
  AN2XD1BWP U673 ( .A1(cu0_RegisterBlock_io_passDataOut_2[3]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4403) );
  AN2XD1BWP U674 ( .A1(cu0_RegisterBlock_io_passDataOut_2[5]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4397) );
  AN2XD1BWP U675 ( .A1(cu0_RegisterBlock_io_passDataOut_2[6]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4394) );
  AN2XD1BWP U676 ( .A1(cu0_RegisterBlock_io_passDataOut_3[0]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4412) );
  AN2XD1BWP U677 ( .A1(cu0_RegisterBlock_io_passDataOut_2[2]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4406) );
  AN2XD1BWP U678 ( .A1(cu0_RegisterBlock_io_passDataOut_2[1]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_4_net4409) );
  AN2XD1BWP U679 ( .A1(cu0_RegisterBlock_io_passDataOut_3[4]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4400) );
  AN2XD1BWP U680 ( .A1(cu0_RegisterBlock_io_passDataOut_3[2]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4406) );
  AN2XD1BWP U681 ( .A1(cu0_RegisterBlock_io_passDataOut_3[6]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4394) );
  AN2XD1BWP U682 ( .A1(cu0_RegisterBlock_io_passDataOut_3[3]), .A2(n333), .Z(
        cu0_RegisterBlock_1_FF_5_net4403) );
  INR2D1BWP U683 ( .A1(cu1_RegisterBlock_FF_io_data_out_6_), .B1(n268), .ZN(
        n267) );
  AN2D1BWP U684 ( .A1(cu1_RegisterBlock_1_FF_1_io_data_out_7_), .A2(n268), .Z(
        n271) );
  CKND2BWP U685 ( .I(cu1_IntFU_1_m_T3[7]), .ZN(n272) );
  NR2D2BWP U686 ( .A1(n272), .A2(n332), .ZN(cu1_RegisterBlock_1_FF_1_net4391)
         );
  CKAN2D1BWP U687 ( .A1(cu0_mem0_io_rdata_0_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4412) );
  CKAN2D1BWP U688 ( .A1(cu0_mem0_io_rdata_1_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4409) );
  CKAN2D1BWP U689 ( .A1(io_command), .A2(n333), .Z(controlBox_N6) );
  CKAN2D1BWP U690 ( .A1(cu0_mem0_io_rdata_3_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4403) );
  CKAN2D1BWP U691 ( .A1(cu0_mem0_io_rdata_4_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4400) );
  CKAN2D1BWP U692 ( .A1(cu0_mem0_io_rdata_2_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4406) );
  CKAN2D1BWP U693 ( .A1(cu0_mem0_io_rdata_6_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4394) );
  CKAN2D1BWP U694 ( .A1(cu0_mem0_io_rdata_7_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4391) );
  CKAN2D1BWP U695 ( .A1(cu0_mem1_io_rdata_0_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4412) );
  CKAN2D1BWP U696 ( .A1(cu0_mem1_io_rdata_1_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4409) );
  CKAN2D1BWP U697 ( .A1(cu0_mem1_io_rdata_2_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4406) );
  CKAN2D1BWP U698 ( .A1(cu0_mem1_io_rdata_3_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4403) );
  CKAN2D1BWP U699 ( .A1(cu0_mem1_io_rdata_4_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4400) );
  CKAN2D1BWP U700 ( .A1(cu0_mem1_io_rdata_5_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4397) );
  CKAN2D1BWP U701 ( .A1(cu0_mem1_io_rdata_6_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4394) );
  CKAN2D1BWP U702 ( .A1(cu0_mem1_io_rdata_7_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_5_net4391) );
  CKAN2D1BWP U703 ( .A1(cu1_mem0_io_rdata_0_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4412) );
  CKAN2D1BWP U704 ( .A1(cu1_mem0_io_rdata_1_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4409) );
  CKAN2D1BWP U705 ( .A1(cu1_mem0_io_rdata_2_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4406) );
  CKAN2D1BWP U706 ( .A1(cu1_mem0_io_rdata_4_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4400) );
  CKAN2D1BWP U707 ( .A1(cu1_mem0_io_rdata_5_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4397) );
  CKAN2D1BWP U708 ( .A1(cu1_mem0_io_rdata_6_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4394) );
  CKAN2D1BWP U709 ( .A1(cu1_mem0_io_rdata_7_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4391) );
  CKAN2D1BWP U710 ( .A1(cu1_mem1_io_rdata_0_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4412) );
  CKAN2D1BWP U711 ( .A1(cu0_mem0_io_rdata_5_), .A2(n333), .Z(
        cu0_RegisterBlock_FF_4_net4397) );
  CKAN2D1BWP U712 ( .A1(cu1_mem1_io_rdata_1_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4409) );
  CKAN2D1BWP U713 ( .A1(cu1_mem1_io_rdata_2_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4406) );
  CKAN2D1BWP U714 ( .A1(cu1_mem1_io_rdata_3_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4403) );
  CKAN2D1BWP U715 ( .A1(cu1_mem1_io_rdata_4_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4400) );
  CKAN2D1BWP U716 ( .A1(cu1_mem1_io_rdata_5_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4397) );
  CKAN2D1BWP U717 ( .A1(cu1_mem1_io_rdata_6_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4394) );
  CKAN2D1BWP U718 ( .A1(cu1_mem0_io_rdata_3_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_4_net4403) );
  CKAN2D1BWP U719 ( .A1(cu1_mem1_io_rdata_7_), .A2(n333), .Z(
        cu1_RegisterBlock_FF_5_net4391) );
  CKND1BWP U720 ( .I(cu0_counterChain_io_data_0_out_2_), .ZN(n275) );
  NR2D1BWP U721 ( .A1(n275), .A2(n332), .ZN(cu0_RegisterBlock_FF_2_net4406) );
  XNR2D1BWP U722 ( .A1(cu0_counterChain_io_data_1_out_0_), .A2(
        cu0_counterChain_io_data_1_out_1_), .ZN(n273) );
  NR2D1BWP U723 ( .A1(n273), .A2(n326), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net4409) );
  XNR2D1BWP U724 ( .A1(cu1_counterChain_io_data_1_out_0_), .A2(
        cu1_counterChain_io_data_1_out_1_), .ZN(n274) );
  NR2D1BWP U725 ( .A1(n274), .A2(n330), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net4409) );
  XNR2D1BWP U726 ( .A1(cu0_counterChain_io_data_0_out_0_), .A2(
        cu0_counterChain_io_data_0_out_1_), .ZN(n276) );
  ND3D1BWP U727 ( .A1(n275), .A2(n333), .A3(
        cu1_counterChain_CounterRC_config__stride_0_), .ZN(n324) );
  NR2D1BWP U728 ( .A1(n276), .A2(n324), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net4409) );
  XNR2D1BWP U729 ( .A1(cu1_counterChain_io_data_0_out_0_), .A2(
        cu1_counterChain_io_data_0_out_1_), .ZN(n277) );
  NR2D1BWP U730 ( .A1(n277), .A2(n328), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net4409) );
  AO22D1BWP U731 ( .A1(n278), .A2(n285), .B1(n298), .B2(
        cu0_counterChain_io_data_1_out_0_), .Z(cu0_RegisterBlock_FF_3_net4412)
         );
  AO22D1BWP U732 ( .A1(n279), .A2(n285), .B1(n298), .B2(
        cu1_counterChain_io_data_1_out_0_), .Z(cu1_RegisterBlock_FF_3_net4412)
         );
  CKND1BWP U733 ( .I(cu0_mem1raMux_io_out_0[0]), .ZN(n280) );
  NR2D1BWP U734 ( .A1(reset), .A2(n280), .ZN(cu0_RegisterBlock_FF_1_net4412)
         );
  AO22D1BWP U735 ( .A1(n281), .A2(n285), .B1(n298), .B2(
        cu0_counterChain_io_data_1_out_1_), .Z(cu0_RegisterBlock_FF_3_net4409)
         );
  AO22D1BWP U736 ( .A1(n282), .A2(n285), .B1(n298), .B2(
        cu1_counterChain_io_data_1_out_1_), .Z(cu1_RegisterBlock_FF_3_net4409)
         );
  AO22D1BWP U737 ( .A1(n283), .A2(n285), .B1(n298), .B2(
        cu1_counterChain_io_data_1_out_2_), .Z(cu1_RegisterBlock_FF_3_net4406)
         );
  AO22D1BWP U738 ( .A1(n284), .A2(n285), .B1(n298), .B2(
        cu0_counterChain_io_data_1_out_2_), .Z(cu0_RegisterBlock_FF_3_net4406)
         );
  CKND1BWP U739 ( .I(n285), .ZN(n289) );
  CKND1BWP U740 ( .I(cu1_mem0raMux_io_out_0[2]), .ZN(n287) );
  NR2D1BWP U741 ( .A1(reset), .A2(n287), .ZN(cu1_RegisterBlock_FF_1_net4406)
         );
  IOA21D1BWP U742 ( .A1(n293), .A2(n298), .B(n292), .ZN(
        cu0_RegisterBlock_FF_1_net4400) );
  IND2D1BWP U744 ( .A1(io_config_enable), .B1(n333), .ZN(
        cu0_controlBlock_incXbar_net4496) );
  NR2D1BWP U745 ( .A1(n299), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_3_net4409)
         );
  NR2D1BWP U746 ( .A1(n300), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_3_net4406)
         );
  NR2D1BWP U747 ( .A1(n301), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_3_net4403)
         );
  NR2D1BWP U748 ( .A1(n302), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_3_net4400)
         );
  NR2D1BWP U749 ( .A1(n303), .A2(reset), .ZN(cu0_RegisterBlock_1_FF_3_net4397)
         );
  NR2D1BWP U750 ( .A1(reset), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net4478) );
  INR2D1BWP U751 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__net4478), .B1(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n304) );
  AO31D1BWP U752 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n333), .B(n304), 
        .Z(cu1_controlBlock_UpDownCtr_1_reg__net4475) );
  NR2D1BWP U753 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n306) );
  CKND1BWP U754 ( .I(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n305) );
  ND2D1BWP U755 ( .A1(n304), .A2(n305), .ZN(n308) );
  OAI31D1BWP U756 ( .A1(reset), .A2(n306), .A3(n305), .B(n308), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net4472) );
  OAI31D1BWP U757 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n307) );
  OAI22D1BWP U758 ( .A1(cu1_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n308), .B1(reset), .B2(n307), .ZN(
        cu1_controlBlock_UpDownCtr_1_reg__net4469) );
  NR2D1BWP U759 ( .A1(reset), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net4478) );
  INR2D1BWP U760 ( .A1(cu0_controlBlock_UpDownCtr_reg__net4478), .B1(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n309) );
  AO31D1BWP U761 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n333), .B(n309), 
        .Z(cu0_controlBlock_UpDownCtr_reg__net4475) );
  NR2D1BWP U762 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n311) );
  CKND1BWP U763 ( .I(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(n310) );
  ND2D1BWP U764 ( .A1(n309), .A2(n310), .ZN(n313) );
  OAI31D1BWP U765 ( .A1(reset), .A2(n311), .A3(n310), .B(n313), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net4472) );
  OAI31D1BWP U766 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n312) );
  OAI22D1BWP U767 ( .A1(cu0_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n313), .B1(reset), .B2(n312), .ZN(
        cu0_controlBlock_UpDownCtr_reg__net4469) );
  NR2D1BWP U768 ( .A1(reset), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net4478) );
  INR2D1BWP U769 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__net4478), .B1(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n314) );
  AO31D1BWP U770 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .A3(n333), .B(n314), 
        .Z(cu0_controlBlock_UpDownCtr_1_reg__net4475) );
  NR2D1BWP U771 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A2(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .ZN(n316) );
  CKND1BWP U772 ( .I(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), .ZN(
        n315) );
  ND2D1BWP U773 ( .A1(n314), .A2(n315), .ZN(n318) );
  OAI31D1BWP U774 ( .A1(reset), .A2(n316), .A3(n315), .B(n318), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net4472) );
  OAI31D1BWP U775 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_2_), 
        .A2(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_0_), .A3(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_1_), .B(
        cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), .ZN(n317) );
  OAI22D1BWP U776 ( .A1(cu0_controlBlock_UpDownCtr_1_reg__io_data_out_3_), 
        .A2(n318), .B1(reset), .B2(n317), .ZN(
        cu0_controlBlock_UpDownCtr_1_reg__net4469) );
  NR2D1BWP U777 ( .A1(reset), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net4478) );
  INR2D1BWP U778 ( .A1(cu1_controlBlock_UpDownCtr_reg__net4478), .B1(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n319) );
  AO31D1BWP U779 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .A3(n333), .B(n319), 
        .Z(cu1_controlBlock_UpDownCtr_reg__net4475) );
  NR2D1BWP U780 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .ZN(n321) );
  CKND1BWP U781 ( .I(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .ZN(n320) );
  ND2D1BWP U782 ( .A1(n319), .A2(n320), .ZN(n323) );
  OAI31D1BWP U783 ( .A1(reset), .A2(n321), .A3(n320), .B(n323), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net4472) );
  OAI31D1BWP U784 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_2_), .A2(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_0_), .A3(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_1_), .B(
        cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .ZN(n322) );
  OAI22D1BWP U785 ( .A1(cu1_controlBlock_UpDownCtr_reg__io_data_out_3_), .A2(
        n323), .B1(reset), .B2(n322), .ZN(
        cu1_controlBlock_UpDownCtr_reg__net4469) );
  NR2D1BWP U786 ( .A1(n324), .A2(cu0_counterChain_io_data_0_out_0_), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net4412) );
  CKND2D1BWP U787 ( .A1(cu0_counterChain_io_data_0_out_0_), .A2(
        cu0_counterChain_io_data_0_out_1_), .ZN(n325) );
  NR2D1BWP U788 ( .A1(n325), .A2(n324), .ZN(
        cu0_counterChain_CounterRC_counter_reg__net4406) );
  NR2D1BWP U789 ( .A1(n326), .A2(cu0_counterChain_io_data_1_out_0_), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net4412) );
  CKND2D1BWP U790 ( .A1(cu0_counterChain_io_data_1_out_0_), .A2(
        cu0_counterChain_io_data_1_out_1_), .ZN(n327) );
  NR2D1BWP U791 ( .A1(n327), .A2(n326), .ZN(
        cu0_counterChain_CounterRC_1_counter_reg__net4406) );
  NR2D1BWP U792 ( .A1(n328), .A2(cu1_counterChain_io_data_0_out_0_), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net4412) );
  CKND2D1BWP U793 ( .A1(cu1_counterChain_io_data_0_out_0_), .A2(
        cu1_counterChain_io_data_0_out_1_), .ZN(n329) );
  NR2D1BWP U794 ( .A1(n329), .A2(n328), .ZN(
        cu1_counterChain_CounterRC_counter_reg__net4406) );
  NR2D1BWP U795 ( .A1(n330), .A2(cu1_counterChain_io_data_1_out_0_), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net4412) );
  CKND2D1BWP U796 ( .A1(cu1_counterChain_io_data_1_out_0_), .A2(
        cu1_counterChain_io_data_1_out_1_), .ZN(n331) );
  NR2D1BWP U797 ( .A1(n331), .A2(n330), .ZN(
        cu1_counterChain_CounterRC_1_counter_reg__net4406) );
endmodule

